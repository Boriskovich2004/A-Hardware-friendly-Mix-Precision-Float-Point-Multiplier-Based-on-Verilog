
module top ( clk, rst_n, data_type, enter, ce, in1_row, in1_col, in2_row, 
        in2_col, disp1_seg, disp1_sel, disp2_seg, disp2_sel, out_seg, out_sel, 
        ready, overflow, error );
  input [3:0] in1_row;
  input [3:0] in1_col;
  input [3:0] in2_row;
  input [3:0] in2_col;
  output [6:0] disp1_seg;
  output [7:0] disp1_sel;
  output [6:0] disp2_seg;
  output [7:0] disp2_sel;
  output [6:0] out_seg;
  output [7:0] out_sel;
  input clk, rst_n, data_type, enter, ce;
  output ready, overflow, error;
  wire   n5007, N1420, N1421, N1422, N1423, N1424, N1425, N1426, N1427, N1428,
         N1429, N1430, N1431, N1432, N1433, N1434, N1435, N1436, N1437, N1438,
         N1439, N1440, N1441, N1442, N1443, N1444, N1445, N1446, N1447, N1448,
         N1449, N1450, N1451, N2679, N2680, N2681, N2682, N2683, N2684, N2685,
         N2686, N2687, N2688, N2689, N2690, N2691, N2692, N2693, N2694, N2695,
         N2696, N2697, N2698, N2699, N2700, N2701, N2702, N2703, N2704, N2705,
         N2706, N2707, N2708, N2709, N2710, N2785, N2786, N2787, N2788, N2789,
         N2790, N2791, N2864, N2865, N2866, N2867, N2868, N2869, N2870, N2943,
         N2944, N2945, N2946, N2947, N2948, N2949, N3022, N3023, N3024, N3025,
         N3026, N3027, N3028, N3172, N3173, N3174, N3175, N3176, N3177, N3178,
         N3324, N3325, N3326, N3327, N3328, N3329, N3330, N3476, N3477, N3478,
         N3479, N3480, N3481, N3482, N3628, N3629, N3630, N3631, N3632, N3633,
         N3634, N3709, N3710, N3711, N3712, N3713, N3714, N3715, N3788, N3789,
         N3790, N3791, N3792, N3793, N3794, N3867, N3868, N3869, N3870, N3871,
         N3872, N3873, N3946, N3947, N3948, N3949, N3950, N3951, N3952, N4096,
         N4097, N4098, N4099, N4100, N4101, N4102, N4248, N4249, N4250, N4251,
         N4252, N4253, N4254, N4400, N4401, N4402, N4403, N4404, N4405, N4406,
         N4552, N4553, N4554, N4555, N4556, N4557, N4558, N4616, N4617, N4618,
         N4619, N4620, N4621, N4622, N4678, N4679, N4680, N4681, N4682, N4683,
         N4684, N4740, N4741, N4742, N4743, N4744, N4745, N4746, N4802, N4803,
         N4804, N4805, N4806, N4807, N4808, N4916, N4917, N4918, N4919, N4920,
         N4921, N4922, N5030, N5031, N5032, N5033, N5034, N5035, N5036, N5144,
         N5145, N5146, N5147, N5148, N5149, N5150, N5258, N5259, N5260, N5261,
         N5262, N5263, N5264, N5268, N5269, N5271, N5294, N5320, N5321, N5323,
         N5346, N5398, \uut/mant_out[0] , \uut/mant_out[1] , \uut/mant_out[2] ,
         \uut/mant_out[3] , \uut/mant_out[4] , \uut/mant_out[5] ,
         \uut/mant_out[6] , \uut/mant_out[7] , \uut/mant_out[8] ,
         \uut/mant_out[9] , \uut/mant_out[10] , \uut/mant_out[11] ,
         \uut/mant_out[12] , \uut/mant_out[13] , \uut/mant_out[14] ,
         \uut/mant_out[15] , \uut/mant_out[16] , \uut/mant_out[17] ,
         \uut/mant_out[18] , \uut/mant_out[19] , \uut/mant_out[20] ,
         \uut/mant_out[21] , \uut/mant_out[22] , \uut/N66 , \uut/start ,
         \uut/N64 , \uut/mult_ready , \uut/normalize , \uut/exp_complete ,
         \uut/valid_q , \uut/more_than_1 , \uut/exp_out[0] , \uut/exp_out[1] ,
         \uut/exp_out[2] , \uut/exp_out[3] , \uut/exp_out[4] ,
         \uut/exp_out[5] , \uut/exp_out[6] , \uut/exp_out[7] ,
         \uut/exp_out[8] , \uut/in2_16_reg[0] , \uut/in2_16_reg[1] ,
         \uut/in2_16_reg[2] , \uut/in2_16_reg[3] , \uut/in2_16_reg[4] ,
         \uut/in2_16_reg[5] , \uut/in2_16_reg[6] , \uut/in2_16_reg[7] ,
         \uut/in2_16_reg[8] , \uut/in2_16_reg[9] , \uut/in2_16_reg[10] ,
         \uut/in2_16_reg[11] , \uut/in2_16_reg[12] , \uut/in2_16_reg[13] ,
         \uut/in2_16_reg[14] , \uut/in2_16_reg[15] , \uut/in1_16_reg[0] ,
         \uut/in1_16_reg[1] , \uut/in1_16_reg[2] , \uut/in1_16_reg[3] ,
         \uut/in1_16_reg[4] , \uut/in1_16_reg[5] , \uut/in1_16_reg[6] ,
         \uut/in1_16_reg[7] , \uut/in1_16_reg[8] , \uut/in1_16_reg[9] ,
         \uut/in1_16_reg[10] , \uut/in1_16_reg[11] , \uut/in1_16_reg[12] ,
         \uut/in1_16_reg[13] , \uut/in1_16_reg[14] , \uut/in1_16_reg[15] ,
         \uut/in2_32_reg[0] , \uut/in2_32_reg[1] , \uut/in2_32_reg[2] ,
         \uut/in2_32_reg[3] , \uut/in2_32_reg[4] , \uut/in2_32_reg[5] ,
         \uut/in2_32_reg[6] , \uut/in2_32_reg[7] , \uut/in2_32_reg[8] ,
         \uut/in2_32_reg[9] , \uut/in2_32_reg[10] , \uut/in2_32_reg[11] ,
         \uut/in2_32_reg[12] , \uut/in2_32_reg[13] , \uut/in2_32_reg[14] ,
         \uut/in2_32_reg[15] , \uut/in2_32_reg[16] , \uut/in2_32_reg[17] ,
         \uut/in2_32_reg[18] , \uut/in2_32_reg[19] , \uut/in2_32_reg[20] ,
         \uut/in2_32_reg[21] , \uut/in2_32_reg[22] , \uut/in2_32_reg[23] ,
         \uut/in2_32_reg[24] , \uut/in2_32_reg[25] , \uut/in2_32_reg[26] ,
         \uut/in2_32_reg[27] , \uut/in2_32_reg[28] , \uut/in2_32_reg[29] ,
         \uut/in2_32_reg[30] , \uut/in2_32_reg[31] , \uut/in1_32_reg[0] ,
         \uut/in1_32_reg[1] , \uut/in1_32_reg[2] , \uut/in1_32_reg[3] ,
         \uut/in1_32_reg[4] , \uut/in1_32_reg[5] , \uut/in1_32_reg[6] ,
         \uut/in1_32_reg[7] , \uut/in1_32_reg[8] , \uut/in1_32_reg[9] ,
         \uut/in1_32_reg[10] , \uut/in1_32_reg[11] , \uut/in1_32_reg[12] ,
         \uut/in1_32_reg[13] , \uut/in1_32_reg[14] , \uut/in1_32_reg[15] ,
         \uut/in1_32_reg[16] , \uut/in1_32_reg[17] , \uut/in1_32_reg[18] ,
         \uut/in1_32_reg[19] , \uut/in1_32_reg[20] , \uut/in1_32_reg[21] ,
         \uut/in1_32_reg[22] , \uut/in1_32_reg[23] , \uut/in1_32_reg[24] ,
         \uut/in1_32_reg[25] , \uut/in1_32_reg[26] , \uut/in1_32_reg[27] ,
         \uut/in1_32_reg[28] , \uut/in1_32_reg[29] , \uut/in1_32_reg[30] ,
         \uut/in1_32_reg[31] , \uut/mult_mant/N299 , \uut/mult_mant/N298 ,
         \uut/mult_mant/temp_product[0] , \uut/mult_mant/temp_product[1] ,
         \uut/mult_mant/temp_product[2] , \uut/mult_mant/temp_product[3] ,
         \uut/mult_mant/temp_product[4] , \uut/mult_mant/temp_product[5] ,
         \uut/mult_mant/temp_product[6] , \uut/mult_mant/temp_product[7] ,
         \uut/mult_mant/temp_product[8] , \uut/mult_mant/temp_product[9] ,
         \uut/mult_mant/temp_product[10] , \uut/mult_mant/temp_product[11] ,
         \uut/mult_mant/temp_product[12] , \uut/mult_mant/temp_product[13] ,
         \uut/mult_mant/temp_product[14] , \uut/mult_mant/temp_product[15] ,
         \uut/mult_mant/temp_product[16] , \uut/mult_mant/temp_product[17] ,
         \uut/mult_mant/temp_product[18] , \uut/mult_mant/temp_product[19] ,
         \uut/mult_mant/temp_product[20] , \uut/mult_mant/temp_product[21] ,
         \uut/mult_mant/temp_product[22] , \uut/mult_mant/temp_product[23] ,
         \uut/mult_mant/temp_product[24] , \uut/mult_mant/temp_product[25] ,
         \uut/mult_mant/temp_product[26] , \uut/mult_mant/temp_product[27] ,
         \uut/mult_mant/temp_product[28] , \uut/mult_mant/temp_product[29] ,
         \uut/mult_mant/temp_product[30] , \uut/mult_mant/temp_product[31] ,
         \uut/mult_mant/temp_product[32] , \uut/mult_mant/temp_product[33] ,
         \uut/mult_mant/temp_product[34] , \uut/mult_mant/temp_product[35] ,
         \uut/mult_mant/temp_product[36] , \uut/mult_mant/temp_product[37] ,
         \uut/mult_mant/temp_product[38] , \uut/mult_mant/temp_product[39] ,
         \uut/mult_mant/temp_product[40] , \uut/mult_mant/temp_product[41] ,
         \uut/mult_mant/temp_product[42] , \uut/mult_mant/temp_product[43] ,
         \uut/mult_mant/temp_product[44] , \uut/mult_mant/temp_product[45] ,
         \uut/mult_mant/temp_product[46] , \uut/mult_mant/temp_product[47] ,
         \uut/mult_mant/mult8_cnt[0] , \uut/mult_mant/mult8_cnt[1] ,
         \uut/mult_mant/mult8_cnt[2] , \uut/mult_mant/mult8_cnt[3] ,
         \uut/mult_mant/state[0] , \uut/mult_mant/state[1] ,
         \uut/mult_mant/state[2] , n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2487, n2488, n2489, n2491, n2493, n2494,
         n2495, n2497, n4991, n4990, n4989, n4994, n4993, n4992, n4997, n4996,
         n4995, n5000, n4999, n4998, n5003, n5002, n5001, n5006, n5005, n5004,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2564, n2566, n2568, n2570, n2572,
         n2574, n2576, n2578, n2580, n2582, n2584, n2586, n2588, n2590, n2592,
         n2594, n2596, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2704, n2705, n2707,
         n2709, n2710, n2711, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2724, n2725, n2726, n2727, n2728, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4987, n4988;
  wire   [3:0] in1_row_q;
  wire   [3:0] in1_col_q;
  wire   [3:0] in2_row_q;
  wire   [3:0] in2_col_q;
  wire   [3:0] in1_row_reg;
  wire   [3:0] in1_col_reg;
  wire   [3:0] in2_row_reg;
  wire   [3:0] in2_col_reg;
  wire   [5:0] input1_cnt;
  wire   [5:0] input2_cnt;
  wire   [31:0] in1_disp;
  wire   [31:0] in2_disp;
  wire   [6:0] disp1_bit7;
  wire   [6:0] disp1_bit6;
  wire   [6:0] disp1_bit5;
  wire   [6:0] disp1_bit4;
  wire   [6:0] disp1_bit3;
  wire   [6:0] disp1_bit2;
  wire   [6:0] disp1_bit1;
  wire   [6:0] disp1_bit0;
  wire   [6:0] disp2_bit7;
  wire   [6:0] disp2_bit6;
  wire   [6:0] disp2_bit5;
  wire   [6:0] disp2_bit4;
  wire   [6:0] disp2_bit3;
  wire   [6:0] disp2_bit2;
  wire   [6:0] disp2_bit1;
  wire   [6:0] disp2_bit0;
  wire   [6:0] bit7;
  wire   [6:0] bit6;
  wire   [6:0] bit5;
  wire   [6:0] bit4;
  wire   [6:0] bit3;
  wire   [6:0] bit2;
  wire   [6:0] bit1;
  wire   [6:0] bit0;
  wire   [2:0] disp1_sel_cnt;
  wire   [2:0] disp2_sel_cnt;
  wire   [2:0] out_sel_cnt;
  wire   [5:0] \uut/mult_mant/shift_amount ;
  wire   [3:0] \uut/mult_mant/mult_end ;
  wire   [7:0] \uut/mult_mant/in2_segment ;
  wire   [7:0] \uut/mult_mant/in1_segment ;
  wire   [7:0] \uut/mult_mant/c2 ;
  wire   [7:0] \uut/mult_mant/b2 ;
  wire   [7:0] \uut/mult_mant/a2 ;
  wire   [7:0] \uut/mult_mant/c1 ;
  wire   [7:0] \uut/mult_mant/b1 ;
  wire   [7:0] \uut/mult_mant/a1 ;

  DFFRHQ \in2_row_q_reg[3]  ( .D(in2_row[3]), .CK(clk), .RN(rst_n), .Q(
        in2_row_q[3]) );
  DFFRHQ \in2_row_q_reg[2]  ( .D(in2_row[2]), .CK(clk), .RN(rst_n), .Q(
        in2_row_q[2]) );
  DFFRHQ \in2_row_q_reg[1]  ( .D(in2_row[1]), .CK(clk), .RN(rst_n), .Q(
        in2_row_q[1]) );
  DFFRHQ \in2_row_q_reg[0]  ( .D(in2_row[0]), .CK(clk), .RN(rst_n), .Q(
        in2_row_q[0]) );
  DFFRHQ \in2_col_q_reg[3]  ( .D(in2_col[3]), .CK(clk), .RN(rst_n), .Q(
        in2_col_q[3]) );
  DFFRHQ \in2_col_q_reg[2]  ( .D(in2_col[2]), .CK(clk), .RN(rst_n), .Q(
        in2_col_q[2]) );
  DFFRHQ \in2_col_q_reg[1]  ( .D(in2_col[1]), .CK(clk), .RN(rst_n), .Q(
        in2_col_q[1]) );
  DFFRHQ \in2_col_q_reg[0]  ( .D(in2_col[0]), .CK(clk), .RN(rst_n), .Q(
        in2_col_q[0]) );
  DFFRHQ \in1_row_q_reg[3]  ( .D(in1_row[3]), .CK(clk), .RN(rst_n), .Q(
        in1_row_q[3]) );
  DFFRHQ \in1_row_q_reg[2]  ( .D(in1_row[2]), .CK(clk), .RN(rst_n), .Q(
        in1_row_q[2]) );
  DFFRHQ \in1_row_q_reg[1]  ( .D(in1_row[1]), .CK(clk), .RN(rst_n), .Q(
        in1_row_q[1]) );
  DFFRHQ \in1_row_q_reg[0]  ( .D(in1_row[0]), .CK(clk), .RN(rst_n), .Q(
        in1_row_q[0]) );
  DFFRHQ \in1_col_q_reg[3]  ( .D(in1_col[3]), .CK(clk), .RN(rst_n), .Q(
        in1_col_q[3]) );
  DFFRHQ \in1_col_q_reg[2]  ( .D(in1_col[2]), .CK(clk), .RN(rst_n), .Q(
        in1_col_q[2]) );
  DFFRHQ \in1_col_q_reg[1]  ( .D(in1_col[1]), .CK(clk), .RN(rst_n), .Q(
        in1_col_q[1]) );
  DFFRHQ \in1_col_q_reg[0]  ( .D(in1_col[0]), .CK(clk), .RN(rst_n), .Q(
        in1_col_q[0]) );
  DFFRHQ \in1_row_reg_reg[3]  ( .D(n4962), .CK(clk), .RN(rst_n), .Q(
        in1_row_reg[3]) );
  DFFRHQ \in1_row_reg_reg[2]  ( .D(n4963), .CK(clk), .RN(rst_n), .Q(
        in1_row_reg[2]) );
  DFFRHQ \in1_row_reg_reg[1]  ( .D(n4964), .CK(clk), .RN(rst_n), .Q(
        in1_row_reg[1]) );
  DFFRHQ \in1_row_reg_reg[0]  ( .D(n4965), .CK(clk), .RN(rst_n), .Q(
        in1_row_reg[0]) );
  DFFRHQ \in1_col_reg_reg[3]  ( .D(n4966), .CK(clk), .RN(rst_n), .Q(
        in1_col_reg[3]) );
  DFFRHQ \in1_col_reg_reg[2]  ( .D(n4967), .CK(clk), .RN(rst_n), .Q(
        in1_col_reg[2]) );
  DFFRHQ \in1_col_reg_reg[1]  ( .D(n4968), .CK(clk), .RN(rst_n), .Q(
        in1_col_reg[1]) );
  DFFRHQ \in1_col_reg_reg[0]  ( .D(n4969), .CK(clk), .RN(rst_n), .Q(
        in1_col_reg[0]) );
  DFFRHQ \in2_row_reg_reg[3]  ( .D(n4970), .CK(clk), .RN(rst_n), .Q(
        in2_row_reg[3]) );
  DFFRHQ \in2_row_reg_reg[2]  ( .D(n4971), .CK(clk), .RN(rst_n), .Q(
        in2_row_reg[2]) );
  DFFRHQ \in2_row_reg_reg[1]  ( .D(n4972), .CK(clk), .RN(rst_n), .Q(
        in2_row_reg[1]) );
  DFFRHQ \in2_row_reg_reg[0]  ( .D(n4973), .CK(clk), .RN(rst_n), .Q(
        in2_row_reg[0]) );
  DFFRHQ \in2_col_reg_reg[3]  ( .D(n4974), .CK(clk), .RN(rst_n), .Q(
        in2_col_reg[3]) );
  DFFRHQ \in2_col_reg_reg[2]  ( .D(n4975), .CK(clk), .RN(rst_n), .Q(
        in2_col_reg[2]) );
  DFFRHQ \in2_col_reg_reg[1]  ( .D(n4976), .CK(clk), .RN(rst_n), .Q(
        in2_col_reg[1]) );
  DFFRHQ \in2_col_reg_reg[0]  ( .D(n4977), .CK(clk), .RN(rst_n), .Q(
        in2_col_reg[0]) );
  DFFRHQ \input1_cnt_reg[0]  ( .D(n2497), .CK(clk), .RN(rst_n), .Q(
        input1_cnt[0]) );
  DFFRHQ \input1_cnt_reg[3]  ( .D(n2493), .CK(clk), .RN(rst_n), .Q(
        input1_cnt[3]) );
  DFFRHQ \input1_cnt_reg[2]  ( .D(n2494), .CK(clk), .RN(rst_n), .Q(
        input1_cnt[2]) );
  DFFRHQ \input1_cnt_reg[1]  ( .D(n2495), .CK(clk), .RN(rst_n), .Q(
        input1_cnt[1]) );
  DFFRHQ \input2_cnt_reg[0]  ( .D(n2491), .CK(clk), .RN(rst_n), .Q(
        input2_cnt[0]) );
  DFFRHQ \input2_cnt_reg[3]  ( .D(n2487), .CK(clk), .RN(rst_n), .Q(
        input2_cnt[3]) );
  DFFRHQ \input2_cnt_reg[2]  ( .D(n2488), .CK(clk), .RN(rst_n), .Q(
        input2_cnt[2]) );
  DFFRHQ \input2_cnt_reg[1]  ( .D(n2489), .CK(clk), .RN(rst_n), .Q(
        input2_cnt[1]) );
  DFFRHQ \input1_reg[31]  ( .D(N1451), .CK(clk), .RN(rst_n), .Q(in1_disp[3])
         );
  DFFRHQ \input1_reg[30]  ( .D(N1450), .CK(clk), .RN(rst_n), .Q(in1_disp[2])
         );
  DFFRHQ \input1_reg[29]  ( .D(N1449), .CK(clk), .RN(rst_n), .Q(in1_disp[1])
         );
  DFFRHQ \input1_reg[28]  ( .D(N1448), .CK(clk), .RN(rst_n), .Q(in1_disp[0])
         );
  DFFRHQ \input1_reg[27]  ( .D(N1447), .CK(clk), .RN(rst_n), .Q(in1_disp[7])
         );
  DFFRHQ \input1_reg[26]  ( .D(N1446), .CK(clk), .RN(rst_n), .Q(in1_disp[6])
         );
  DFFRHQ \input1_reg[25]  ( .D(N1445), .CK(clk), .RN(rst_n), .Q(in1_disp[5])
         );
  DFFRHQ \input1_reg[24]  ( .D(N1444), .CK(clk), .RN(rst_n), .Q(in1_disp[4])
         );
  DFFRHQ \input1_reg[23]  ( .D(N1443), .CK(clk), .RN(rst_n), .Q(in1_disp[11])
         );
  DFFRHQ \input1_reg[22]  ( .D(N1442), .CK(clk), .RN(rst_n), .Q(in1_disp[10])
         );
  DFFRHQ \input1_reg[21]  ( .D(N1441), .CK(clk), .RN(rst_n), .Q(in1_disp[9])
         );
  DFFRHQ \input1_reg[20]  ( .D(N1440), .CK(clk), .RN(rst_n), .Q(in1_disp[8])
         );
  DFFRHQ \input1_reg[19]  ( .D(N1439), .CK(clk), .RN(rst_n), .Q(in1_disp[15])
         );
  DFFRHQ \input1_reg[18]  ( .D(N1438), .CK(clk), .RN(rst_n), .Q(in1_disp[14])
         );
  DFFRHQ \input1_reg[17]  ( .D(N1437), .CK(clk), .RN(rst_n), .Q(in1_disp[13])
         );
  DFFRHQ \input1_reg[16]  ( .D(N1436), .CK(clk), .RN(rst_n), .Q(in1_disp[12])
         );
  DFFRHQ \input1_reg[15]  ( .D(N1435), .CK(clk), .RN(rst_n), .Q(in1_disp[19])
         );
  DFFRHQ \input1_reg[14]  ( .D(N1434), .CK(clk), .RN(rst_n), .Q(in1_disp[18])
         );
  DFFRHQ \input1_reg[13]  ( .D(N1433), .CK(clk), .RN(rst_n), .Q(in1_disp[17])
         );
  DFFRHQ \input1_reg[12]  ( .D(N1432), .CK(clk), .RN(rst_n), .Q(in1_disp[16])
         );
  DFFRHQ \input1_reg[11]  ( .D(N1431), .CK(clk), .RN(rst_n), .Q(in1_disp[23])
         );
  DFFRHQ \input1_reg[10]  ( .D(N1430), .CK(clk), .RN(rst_n), .Q(in1_disp[22])
         );
  DFFRHQ \input1_reg[9]  ( .D(N1429), .CK(clk), .RN(rst_n), .Q(in1_disp[21])
         );
  DFFRHQ \input1_reg[8]  ( .D(N1428), .CK(clk), .RN(rst_n), .Q(in1_disp[20])
         );
  DFFRHQ \input1_reg[7]  ( .D(N1427), .CK(clk), .RN(rst_n), .Q(in1_disp[27])
         );
  DFFRHQ \input1_reg[6]  ( .D(N1426), .CK(clk), .RN(rst_n), .Q(in1_disp[26])
         );
  DFFRHQ \input1_reg[5]  ( .D(N1425), .CK(clk), .RN(rst_n), .Q(in1_disp[25])
         );
  DFFRHQ \input1_reg[4]  ( .D(N1424), .CK(clk), .RN(rst_n), .Q(in1_disp[24])
         );
  DFFRHQ \input1_reg[3]  ( .D(N1423), .CK(clk), .RN(rst_n), .Q(in1_disp[31])
         );
  DFFRHQ \input1_reg[2]  ( .D(N1422), .CK(clk), .RN(rst_n), .Q(in1_disp[30])
         );
  DFFRHQ \input1_reg[1]  ( .D(N1421), .CK(clk), .RN(rst_n), .Q(in1_disp[29])
         );
  DFFRHQ \input1_reg[0]  ( .D(N1420), .CK(clk), .RN(rst_n), .Q(in1_disp[28])
         );
  DFFRHQ \input2_reg[31]  ( .D(N2710), .CK(clk), .RN(rst_n), .Q(in2_disp[3])
         );
  DFFRHQ \input2_reg[30]  ( .D(N2709), .CK(clk), .RN(rst_n), .Q(in2_disp[2])
         );
  DFFRHQ \input2_reg[29]  ( .D(N2708), .CK(clk), .RN(rst_n), .Q(in2_disp[1])
         );
  DFFRHQ \input2_reg[28]  ( .D(N2707), .CK(clk), .RN(rst_n), .Q(in2_disp[0])
         );
  DFFRHQ \input2_reg[27]  ( .D(N2706), .CK(clk), .RN(rst_n), .Q(in2_disp[7])
         );
  DFFRHQ \input2_reg[26]  ( .D(N2705), .CK(clk), .RN(rst_n), .Q(in2_disp[6])
         );
  DFFRHQ \input2_reg[25]  ( .D(N2704), .CK(clk), .RN(rst_n), .Q(in2_disp[5])
         );
  DFFRHQ \input2_reg[24]  ( .D(N2703), .CK(clk), .RN(rst_n), .Q(in2_disp[4])
         );
  DFFRHQ \input2_reg[23]  ( .D(N2702), .CK(clk), .RN(rst_n), .Q(in2_disp[11])
         );
  DFFRHQ \input2_reg[22]  ( .D(N2701), .CK(clk), .RN(rst_n), .Q(in2_disp[10])
         );
  DFFRHQ \input2_reg[21]  ( .D(N2700), .CK(clk), .RN(rst_n), .Q(in2_disp[9])
         );
  DFFRHQ \input2_reg[20]  ( .D(N2699), .CK(clk), .RN(rst_n), .Q(in2_disp[8])
         );
  DFFRHQ \input2_reg[19]  ( .D(N2698), .CK(clk), .RN(rst_n), .Q(in2_disp[15])
         );
  DFFRHQ \input2_reg[18]  ( .D(N2697), .CK(clk), .RN(rst_n), .Q(in2_disp[14])
         );
  DFFRHQ \input2_reg[17]  ( .D(N2696), .CK(clk), .RN(rst_n), .Q(in2_disp[13])
         );
  DFFRHQ \input2_reg[16]  ( .D(N2695), .CK(clk), .RN(rst_n), .Q(in2_disp[12])
         );
  DFFRHQ \input2_reg[15]  ( .D(N2694), .CK(clk), .RN(rst_n), .Q(in2_disp[19])
         );
  DFFRHQ \input2_reg[14]  ( .D(N2693), .CK(clk), .RN(rst_n), .Q(in2_disp[18])
         );
  DFFRHQ \input2_reg[13]  ( .D(N2692), .CK(clk), .RN(rst_n), .Q(in2_disp[17])
         );
  DFFRHQ \input2_reg[12]  ( .D(N2691), .CK(clk), .RN(rst_n), .Q(in2_disp[16])
         );
  DFFRHQ \input2_reg[11]  ( .D(N2690), .CK(clk), .RN(rst_n), .Q(in2_disp[23])
         );
  DFFRHQ \input2_reg[10]  ( .D(N2689), .CK(clk), .RN(rst_n), .Q(in2_disp[22])
         );
  DFFRHQ \input2_reg[9]  ( .D(N2688), .CK(clk), .RN(rst_n), .Q(in2_disp[21])
         );
  DFFRHQ \input2_reg[8]  ( .D(N2687), .CK(clk), .RN(rst_n), .Q(in2_disp[20])
         );
  DFFRHQ \input2_reg[7]  ( .D(N2686), .CK(clk), .RN(rst_n), .Q(in2_disp[27])
         );
  DFFRHQ \input2_reg[6]  ( .D(N2685), .CK(clk), .RN(rst_n), .Q(in2_disp[26])
         );
  DFFRHQ \input2_reg[5]  ( .D(N2684), .CK(clk), .RN(rst_n), .Q(in2_disp[25])
         );
  DFFRHQ \input2_reg[4]  ( .D(N2683), .CK(clk), .RN(rst_n), .Q(in2_disp[24])
         );
  DFFRHQ \input2_reg[3]  ( .D(N2682), .CK(clk), .RN(rst_n), .Q(in2_disp[31])
         );
  DFFRHQ \input2_reg[2]  ( .D(N2681), .CK(clk), .RN(rst_n), .Q(in2_disp[30])
         );
  DFFRHQ \input2_reg[1]  ( .D(N2680), .CK(clk), .RN(rst_n), .Q(in2_disp[29])
         );
  DFFRHQ \input2_reg[0]  ( .D(N2679), .CK(clk), .RN(rst_n), .Q(in2_disp[28])
         );
  DFFRHQ \disp1_bit7_reg[6]  ( .D(N2791), .CK(clk), .RN(rst_n), .Q(
        disp1_bit7[6]) );
  DFFRHQ \disp1_bit7_reg[5]  ( .D(N2790), .CK(clk), .RN(rst_n), .Q(
        disp1_bit7[5]) );
  DFFRHQ \disp1_bit7_reg[4]  ( .D(N2789), .CK(clk), .RN(rst_n), .Q(
        disp1_bit7[4]) );
  DFFRHQ \disp1_bit7_reg[3]  ( .D(N2788), .CK(clk), .RN(rst_n), .Q(
        disp1_bit7[3]) );
  DFFRHQ \disp1_bit7_reg[2]  ( .D(N2787), .CK(clk), .RN(rst_n), .Q(
        disp1_bit7[2]) );
  DFFRHQ \disp1_bit7_reg[1]  ( .D(N2786), .CK(clk), .RN(rst_n), .Q(
        disp1_bit7[1]) );
  DFFRHQ \disp1_bit7_reg[0]  ( .D(N2785), .CK(clk), .RN(rst_n), .Q(
        disp1_bit7[0]) );
  DFFRHQ \disp1_bit6_reg[6]  ( .D(N2870), .CK(clk), .RN(rst_n), .Q(
        disp1_bit6[6]) );
  DFFRHQ \disp1_bit6_reg[5]  ( .D(N2869), .CK(clk), .RN(rst_n), .Q(
        disp1_bit6[5]) );
  DFFRHQ \disp1_bit6_reg[4]  ( .D(N2868), .CK(clk), .RN(rst_n), .Q(
        disp1_bit6[4]) );
  DFFRHQ \disp1_bit6_reg[3]  ( .D(N2867), .CK(clk), .RN(rst_n), .Q(
        disp1_bit6[3]) );
  DFFRHQ \disp1_bit6_reg[2]  ( .D(N2866), .CK(clk), .RN(rst_n), .Q(
        disp1_bit6[2]) );
  DFFRHQ \disp1_bit6_reg[1]  ( .D(N2865), .CK(clk), .RN(rst_n), .Q(
        disp1_bit6[1]) );
  DFFRHQ \disp1_bit6_reg[0]  ( .D(N2864), .CK(clk), .RN(rst_n), .Q(
        disp1_bit6[0]) );
  DFFRHQ \disp1_bit5_reg[6]  ( .D(N2949), .CK(clk), .RN(rst_n), .Q(
        disp1_bit5[6]) );
  DFFRHQ \disp1_bit5_reg[5]  ( .D(N2948), .CK(clk), .RN(rst_n), .Q(
        disp1_bit5[5]) );
  DFFRHQ \disp1_bit5_reg[4]  ( .D(N2947), .CK(clk), .RN(rst_n), .Q(
        disp1_bit5[4]) );
  DFFRHQ \disp1_bit5_reg[3]  ( .D(N2946), .CK(clk), .RN(rst_n), .Q(
        disp1_bit5[3]) );
  DFFRHQ \disp1_bit5_reg[2]  ( .D(N2945), .CK(clk), .RN(rst_n), .Q(
        disp1_bit5[2]) );
  DFFRHQ \disp1_bit5_reg[1]  ( .D(N2944), .CK(clk), .RN(rst_n), .Q(
        disp1_bit5[1]) );
  DFFRHQ \disp1_bit5_reg[0]  ( .D(N2943), .CK(clk), .RN(rst_n), .Q(
        disp1_bit5[0]) );
  DFFRHQ \disp1_bit4_reg[6]  ( .D(N3028), .CK(clk), .RN(rst_n), .Q(
        disp1_bit4[6]) );
  DFFRHQ \disp1_bit4_reg[5]  ( .D(N3027), .CK(clk), .RN(rst_n), .Q(
        disp1_bit4[5]) );
  DFFRHQ \disp1_bit4_reg[4]  ( .D(N3026), .CK(clk), .RN(rst_n), .Q(
        disp1_bit4[4]) );
  DFFRHQ \disp1_bit4_reg[3]  ( .D(N3025), .CK(clk), .RN(rst_n), .Q(
        disp1_bit4[3]) );
  DFFRHQ \disp1_bit4_reg[2]  ( .D(N3024), .CK(clk), .RN(rst_n), .Q(
        disp1_bit4[2]) );
  DFFRHQ \disp1_bit4_reg[1]  ( .D(N3023), .CK(clk), .RN(rst_n), .Q(
        disp1_bit4[1]) );
  DFFRHQ \disp1_bit4_reg[0]  ( .D(N3022), .CK(clk), .RN(rst_n), .Q(
        disp1_bit4[0]) );
  DFFRHQ \disp1_bit3_reg[6]  ( .D(N3178), .CK(clk), .RN(rst_n), .Q(
        disp1_bit3[6]) );
  DFFRHQ \disp1_bit3_reg[5]  ( .D(N3177), .CK(clk), .RN(rst_n), .Q(
        disp1_bit3[5]) );
  DFFRHQ \disp1_bit3_reg[4]  ( .D(N3176), .CK(clk), .RN(rst_n), .Q(
        disp1_bit3[4]) );
  DFFRHQ \disp1_bit3_reg[3]  ( .D(N3175), .CK(clk), .RN(rst_n), .Q(
        disp1_bit3[3]) );
  DFFRHQ \disp1_bit3_reg[2]  ( .D(N3174), .CK(clk), .RN(rst_n), .Q(
        disp1_bit3[2]) );
  DFFRHQ \disp1_bit3_reg[1]  ( .D(N3173), .CK(clk), .RN(rst_n), .Q(
        disp1_bit3[1]) );
  DFFRHQ \disp1_bit3_reg[0]  ( .D(N3172), .CK(clk), .RN(rst_n), .Q(
        disp1_bit3[0]) );
  DFFRHQ \disp1_bit2_reg[6]  ( .D(N3330), .CK(clk), .RN(rst_n), .Q(
        disp1_bit2[6]) );
  DFFRHQ \disp1_bit2_reg[5]  ( .D(N3329), .CK(clk), .RN(rst_n), .Q(
        disp1_bit2[5]) );
  DFFRHQ \disp1_bit2_reg[4]  ( .D(N3328), .CK(clk), .RN(rst_n), .Q(
        disp1_bit2[4]) );
  DFFRHQ \disp1_bit2_reg[3]  ( .D(N3327), .CK(clk), .RN(rst_n), .Q(
        disp1_bit2[3]) );
  DFFRHQ \disp1_bit2_reg[2]  ( .D(N3326), .CK(clk), .RN(rst_n), .Q(
        disp1_bit2[2]) );
  DFFRHQ \disp1_bit2_reg[1]  ( .D(N3325), .CK(clk), .RN(rst_n), .Q(
        disp1_bit2[1]) );
  DFFRHQ \disp1_bit2_reg[0]  ( .D(N3324), .CK(clk), .RN(rst_n), .Q(
        disp1_bit2[0]) );
  DFFRHQ \disp1_bit1_reg[6]  ( .D(N3482), .CK(clk), .RN(rst_n), .Q(
        disp1_bit1[6]) );
  DFFRHQ \disp1_bit1_reg[5]  ( .D(N3481), .CK(clk), .RN(rst_n), .Q(
        disp1_bit1[5]) );
  DFFRHQ \disp1_bit1_reg[4]  ( .D(N3480), .CK(clk), .RN(rst_n), .Q(
        disp1_bit1[4]) );
  DFFRHQ \disp1_bit1_reg[3]  ( .D(N3479), .CK(clk), .RN(rst_n), .Q(
        disp1_bit1[3]) );
  DFFRHQ \disp1_bit1_reg[2]  ( .D(N3478), .CK(clk), .RN(rst_n), .Q(
        disp1_bit1[2]) );
  DFFRHQ \disp1_bit1_reg[1]  ( .D(N3477), .CK(clk), .RN(rst_n), .Q(
        disp1_bit1[1]) );
  DFFRHQ \disp1_bit1_reg[0]  ( .D(N3476), .CK(clk), .RN(rst_n), .Q(
        disp1_bit1[0]) );
  DFFRHQ \disp1_bit0_reg[6]  ( .D(N3634), .CK(clk), .RN(rst_n), .Q(
        disp1_bit0[6]) );
  DFFRHQ \disp1_bit0_reg[5]  ( .D(N3633), .CK(clk), .RN(rst_n), .Q(
        disp1_bit0[5]) );
  DFFRHQ \disp1_bit0_reg[4]  ( .D(N3632), .CK(clk), .RN(rst_n), .Q(
        disp1_bit0[4]) );
  DFFRHQ \disp1_bit0_reg[3]  ( .D(N3631), .CK(clk), .RN(rst_n), .Q(
        disp1_bit0[3]) );
  DFFRHQ \disp1_bit0_reg[2]  ( .D(N3630), .CK(clk), .RN(rst_n), .Q(
        disp1_bit0[2]) );
  DFFRHQ \disp1_bit0_reg[1]  ( .D(N3629), .CK(clk), .RN(rst_n), .Q(
        disp1_bit0[1]) );
  DFFRHQ \disp1_bit0_reg[0]  ( .D(N3628), .CK(clk), .RN(rst_n), .Q(
        disp1_bit0[0]) );
  DFFRHQ \disp2_bit7_reg[6]  ( .D(N3715), .CK(clk), .RN(rst_n), .Q(
        disp2_bit7[6]) );
  DFFRHQ \disp2_bit7_reg[5]  ( .D(N3714), .CK(clk), .RN(rst_n), .Q(
        disp2_bit7[5]) );
  DFFRHQ \disp2_bit7_reg[4]  ( .D(N3713), .CK(clk), .RN(rst_n), .Q(
        disp2_bit7[4]) );
  DFFRHQ \disp2_bit7_reg[3]  ( .D(N3712), .CK(clk), .RN(rst_n), .Q(
        disp2_bit7[3]) );
  DFFRHQ \disp2_bit7_reg[2]  ( .D(N3711), .CK(clk), .RN(rst_n), .Q(
        disp2_bit7[2]) );
  DFFRHQ \disp2_bit7_reg[1]  ( .D(N3710), .CK(clk), .RN(rst_n), .Q(
        disp2_bit7[1]) );
  DFFRHQ \disp2_bit7_reg[0]  ( .D(N3709), .CK(clk), .RN(rst_n), .Q(
        disp2_bit7[0]) );
  DFFRHQ \disp2_bit6_reg[6]  ( .D(N3794), .CK(clk), .RN(rst_n), .Q(
        disp2_bit6[6]) );
  DFFRHQ \disp2_bit6_reg[5]  ( .D(N3793), .CK(clk), .RN(rst_n), .Q(
        disp2_bit6[5]) );
  DFFRHQ \disp2_bit6_reg[4]  ( .D(N3792), .CK(clk), .RN(rst_n), .Q(
        disp2_bit6[4]) );
  DFFRHQ \disp2_bit6_reg[3]  ( .D(N3791), .CK(clk), .RN(rst_n), .Q(
        disp2_bit6[3]) );
  DFFRHQ \disp2_bit6_reg[2]  ( .D(N3790), .CK(clk), .RN(rst_n), .Q(
        disp2_bit6[2]) );
  DFFRHQ \disp2_bit6_reg[1]  ( .D(N3789), .CK(clk), .RN(rst_n), .Q(
        disp2_bit6[1]) );
  DFFRHQ \disp2_bit6_reg[0]  ( .D(N3788), .CK(clk), .RN(rst_n), .Q(
        disp2_bit6[0]) );
  DFFRHQ \disp2_bit5_reg[6]  ( .D(N3873), .CK(clk), .RN(rst_n), .Q(
        disp2_bit5[6]) );
  DFFRHQ \disp2_bit5_reg[5]  ( .D(N3872), .CK(clk), .RN(rst_n), .Q(
        disp2_bit5[5]) );
  DFFRHQ \disp2_bit5_reg[4]  ( .D(N3871), .CK(clk), .RN(rst_n), .Q(
        disp2_bit5[4]) );
  DFFRHQ \disp2_bit5_reg[3]  ( .D(N3870), .CK(clk), .RN(rst_n), .Q(
        disp2_bit5[3]) );
  DFFRHQ \disp2_bit5_reg[2]  ( .D(N3869), .CK(clk), .RN(rst_n), .Q(
        disp2_bit5[2]) );
  DFFRHQ \disp2_bit5_reg[1]  ( .D(N3868), .CK(clk), .RN(rst_n), .Q(
        disp2_bit5[1]) );
  DFFRHQ \disp2_bit5_reg[0]  ( .D(N3867), .CK(clk), .RN(rst_n), .Q(
        disp2_bit5[0]) );
  DFFRHQ \disp2_bit4_reg[6]  ( .D(N3952), .CK(clk), .RN(rst_n), .Q(
        disp2_bit4[6]) );
  DFFRHQ \disp2_bit4_reg[5]  ( .D(N3951), .CK(clk), .RN(rst_n), .Q(
        disp2_bit4[5]) );
  DFFRHQ \disp2_bit4_reg[4]  ( .D(N3950), .CK(clk), .RN(rst_n), .Q(
        disp2_bit4[4]) );
  DFFRHQ \disp2_bit4_reg[3]  ( .D(N3949), .CK(clk), .RN(rst_n), .Q(
        disp2_bit4[3]) );
  DFFRHQ \disp2_bit4_reg[2]  ( .D(N3948), .CK(clk), .RN(rst_n), .Q(
        disp2_bit4[2]) );
  DFFRHQ \disp2_bit4_reg[1]  ( .D(N3947), .CK(clk), .RN(rst_n), .Q(
        disp2_bit4[1]) );
  DFFRHQ \disp2_bit4_reg[0]  ( .D(N3946), .CK(clk), .RN(rst_n), .Q(
        disp2_bit4[0]) );
  DFFRHQ \disp2_bit3_reg[6]  ( .D(N4102), .CK(clk), .RN(rst_n), .Q(
        disp2_bit3[6]) );
  DFFRHQ \disp2_bit3_reg[5]  ( .D(N4101), .CK(clk), .RN(rst_n), .Q(
        disp2_bit3[5]) );
  DFFRHQ \disp2_bit3_reg[4]  ( .D(N4100), .CK(clk), .RN(rst_n), .Q(
        disp2_bit3[4]) );
  DFFRHQ \disp2_bit3_reg[3]  ( .D(N4099), .CK(clk), .RN(rst_n), .Q(
        disp2_bit3[3]) );
  DFFRHQ \disp2_bit3_reg[2]  ( .D(N4098), .CK(clk), .RN(rst_n), .Q(
        disp2_bit3[2]) );
  DFFRHQ \disp2_bit3_reg[1]  ( .D(N4097), .CK(clk), .RN(rst_n), .Q(
        disp2_bit3[1]) );
  DFFRHQ \disp2_bit3_reg[0]  ( .D(N4096), .CK(clk), .RN(rst_n), .Q(
        disp2_bit3[0]) );
  DFFRHQ \disp2_bit2_reg[6]  ( .D(N4254), .CK(clk), .RN(rst_n), .Q(
        disp2_bit2[6]) );
  DFFRHQ \disp2_bit2_reg[5]  ( .D(N4253), .CK(clk), .RN(rst_n), .Q(
        disp2_bit2[5]) );
  DFFRHQ \disp2_bit2_reg[4]  ( .D(N4252), .CK(clk), .RN(rst_n), .Q(
        disp2_bit2[4]) );
  DFFRHQ \disp2_bit2_reg[3]  ( .D(N4251), .CK(clk), .RN(rst_n), .Q(
        disp2_bit2[3]) );
  DFFRHQ \disp2_bit2_reg[2]  ( .D(N4250), .CK(clk), .RN(rst_n), .Q(
        disp2_bit2[2]) );
  DFFRHQ \disp2_bit2_reg[1]  ( .D(N4249), .CK(clk), .RN(rst_n), .Q(
        disp2_bit2[1]) );
  DFFRHQ \disp2_bit2_reg[0]  ( .D(N4248), .CK(clk), .RN(rst_n), .Q(
        disp2_bit2[0]) );
  DFFRHQ \disp2_bit1_reg[6]  ( .D(N4406), .CK(clk), .RN(rst_n), .Q(
        disp2_bit1[6]) );
  DFFRHQ \disp2_bit1_reg[5]  ( .D(N4405), .CK(clk), .RN(rst_n), .Q(
        disp2_bit1[5]) );
  DFFRHQ \disp2_bit1_reg[4]  ( .D(N4404), .CK(clk), .RN(rst_n), .Q(
        disp2_bit1[4]) );
  DFFRHQ \disp2_bit1_reg[3]  ( .D(N4403), .CK(clk), .RN(rst_n), .Q(
        disp2_bit1[3]) );
  DFFRHQ \disp2_bit1_reg[2]  ( .D(N4402), .CK(clk), .RN(rst_n), .Q(
        disp2_bit1[2]) );
  DFFRHQ \disp2_bit1_reg[1]  ( .D(N4401), .CK(clk), .RN(rst_n), .Q(
        disp2_bit1[1]) );
  DFFRHQ \disp2_bit1_reg[0]  ( .D(N4400), .CK(clk), .RN(rst_n), .Q(
        disp2_bit1[0]) );
  DFFRHQ \disp2_bit0_reg[6]  ( .D(N4558), .CK(clk), .RN(rst_n), .Q(
        disp2_bit0[6]) );
  DFFRHQ \disp2_bit0_reg[5]  ( .D(N4557), .CK(clk), .RN(rst_n), .Q(
        disp2_bit0[5]) );
  DFFRHQ \disp2_bit0_reg[4]  ( .D(N4556), .CK(clk), .RN(rst_n), .Q(
        disp2_bit0[4]) );
  DFFRHQ \disp2_bit0_reg[3]  ( .D(N4555), .CK(clk), .RN(rst_n), .Q(
        disp2_bit0[3]) );
  DFFRHQ \disp2_bit0_reg[2]  ( .D(N4554), .CK(clk), .RN(rst_n), .Q(
        disp2_bit0[2]) );
  DFFRHQ \disp2_bit0_reg[1]  ( .D(N4553), .CK(clk), .RN(rst_n), .Q(
        disp2_bit0[1]) );
  DFFRHQ \disp2_bit0_reg[0]  ( .D(N4552), .CK(clk), .RN(rst_n), .Q(
        disp2_bit0[0]) );
  DFFRHQ \disp1_sel_cnt_reg[0]  ( .D(n4978), .CK(clk), .RN(rst_n), .Q(
        disp1_sel_cnt[0]) );
  DFFRHQ \disp1_sel_cnt_reg[1]  ( .D(N5268), .CK(clk), .RN(rst_n), .Q(
        disp1_sel_cnt[1]) );
  DFFRHQ \disp1_sel_cnt_reg[2]  ( .D(N5269), .CK(clk), .RN(rst_n), .Q(
        disp1_sel_cnt[2]) );
  DFFRHQ \disp2_sel_cnt_reg[0]  ( .D(n4979), .CK(clk), .RN(rst_n), .Q(
        disp2_sel_cnt[0]) );
  DFFRHQ \disp2_sel_cnt_reg[1]  ( .D(N5320), .CK(clk), .RN(rst_n), .Q(
        disp2_sel_cnt[1]) );
  DFFRHQ \disp2_sel_cnt_reg[2]  ( .D(N5321), .CK(clk), .RN(rst_n), .Q(
        disp2_sel_cnt[2]) );
  DFFRHQ \out_sel_cnt_reg[2]  ( .D(N5321), .CK(clk), .RN(rst_n), .Q(
        out_sel_cnt[2]) );
  DFFRHQ \out_sel_cnt_reg[1]  ( .D(N5320), .CK(clk), .RN(rst_n), .Q(
        out_sel_cnt[1]) );
  DFFRHQ \out_sel_cnt_reg[0]  ( .D(n4979), .CK(clk), .RN(rst_n), .Q(
        out_sel_cnt[0]) );
  DFFRHQ \uut/valid_q_reg  ( .D(enter), .CK(clk), .RN(rst_n), .Q(\uut/valid_q ) );
  DFFRHQ \uut/mult_mant/mult_end_reg[2]  ( .D(n4961), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/mult_end [2]) );
  DFFRHQ \uut/mult_mant/mult_end_reg[3]  ( .D(data_type), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/mult_end [3]) );
  DFFRHQ \uut/mult_mant/state_reg[0]  ( .D(\uut/mult_mant/N298 ), .CK(clk), 
        .RN(rst_n), .Q(\uut/mult_mant/state[0] ) );
  DFFRHQ \uut/mult_mant/state_reg[1]  ( .D(\uut/mult_mant/N299 ), .CK(clk), 
        .RN(rst_n), .Q(\uut/mult_mant/state[1] ) );
  DFFRHQ \uut/mult_mant/state_reg[2]  ( .D(n2641), .CK(clk), .RN(rst_n), .Q(
        \uut/mult_mant/state[2] ) );
  DFFSHQ \uut/mult_mant/ready_reg  ( .D(n2485), .CK(clk), .SN(rst_n), .Q(
        \uut/mult_ready ) );
  DFFSHQ \uut/ready_reg  ( .D(\uut/N64 ), .CK(clk), .SN(rst_n), .Q(ready) );
  DFFRHQ \uut/in1_32_reg_reg[31]  ( .D(n2400), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[31] ) );
  DFFRHQ \uut/in1_32_reg_reg[30]  ( .D(n2399), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[30] ) );
  DFFRHQ \uut/in1_32_reg_reg[29]  ( .D(n2398), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[29] ) );
  DFFRHQ \uut/in1_32_reg_reg[28]  ( .D(n2397), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[28] ) );
  DFFRHQ \uut/in1_32_reg_reg[27]  ( .D(n2396), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[27] ) );
  DFFRHQ \uut/in1_32_reg_reg[26]  ( .D(n2395), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[26] ) );
  DFFRHQ \uut/in1_32_reg_reg[25]  ( .D(n2394), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[25] ) );
  DFFRHQ \uut/in1_32_reg_reg[24]  ( .D(n2393), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[24] ) );
  DFFRHQ \uut/in1_32_reg_reg[23]  ( .D(n2392), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[23] ) );
  DFFRHQ \uut/in1_32_reg_reg[22]  ( .D(n2391), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[22] ) );
  DFFRHQ \uut/in1_32_reg_reg[21]  ( .D(n2390), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[21] ) );
  DFFRHQ \uut/in1_32_reg_reg[20]  ( .D(n2389), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[20] ) );
  DFFRHQ \uut/in1_32_reg_reg[19]  ( .D(n2388), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[19] ) );
  DFFRHQ \uut/in1_32_reg_reg[18]  ( .D(n2387), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[18] ) );
  DFFRHQ \uut/in1_32_reg_reg[17]  ( .D(n2386), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[17] ) );
  DFFRHQ \uut/in1_32_reg_reg[16]  ( .D(n2385), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[16] ) );
  DFFRHQ \uut/in1_32_reg_reg[15]  ( .D(n2384), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[15] ) );
  DFFRHQ \uut/in1_32_reg_reg[14]  ( .D(n2383), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[14] ) );
  DFFRHQ \uut/in1_32_reg_reg[13]  ( .D(n2382), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[13] ) );
  DFFRHQ \uut/in1_32_reg_reg[12]  ( .D(n2381), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[12] ) );
  DFFRHQ \uut/in1_32_reg_reg[11]  ( .D(n2380), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[11] ) );
  DFFRHQ \uut/in1_32_reg_reg[10]  ( .D(n2379), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[10] ) );
  DFFRHQ \uut/in1_32_reg_reg[9]  ( .D(n2378), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[9] ) );
  DFFRHQ \uut/in1_32_reg_reg[8]  ( .D(n2377), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[8] ) );
  DFFRHQ \uut/in1_32_reg_reg[7]  ( .D(n2376), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[7] ) );
  DFFRHQ \uut/in1_32_reg_reg[6]  ( .D(n2375), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[6] ) );
  DFFRHQ \uut/in1_32_reg_reg[5]  ( .D(n2374), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[5] ) );
  DFFRHQ \uut/in1_32_reg_reg[4]  ( .D(n2373), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[4] ) );
  DFFRHQ \uut/in1_32_reg_reg[3]  ( .D(n2372), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[3] ) );
  DFFRHQ \uut/in1_32_reg_reg[2]  ( .D(n2371), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[2] ) );
  DFFRHQ \uut/in1_32_reg_reg[1]  ( .D(n2370), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[1] ) );
  DFFRHQ \uut/in1_32_reg_reg[0]  ( .D(n2369), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_32_reg[0] ) );
  DFFRHQ \uut/in2_32_reg_reg[31]  ( .D(n2368), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[31] ) );
  DFFRHQ \uut/in2_32_reg_reg[30]  ( .D(n2367), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[30] ) );
  DFFRHQ \uut/in2_32_reg_reg[29]  ( .D(n2366), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[29] ) );
  DFFRHQ \uut/in2_32_reg_reg[28]  ( .D(n2365), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[28] ) );
  DFFRHQ \uut/in2_32_reg_reg[27]  ( .D(n2364), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[27] ) );
  DFFRHQ \uut/in2_32_reg_reg[26]  ( .D(n2363), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[26] ) );
  DFFRHQ \uut/in2_32_reg_reg[25]  ( .D(n2362), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[25] ) );
  DFFRHQ \uut/in2_32_reg_reg[24]  ( .D(n2361), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[24] ) );
  DFFRHQ \uut/in2_32_reg_reg[23]  ( .D(n2360), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[23] ) );
  DFFRHQ \uut/in2_32_reg_reg[22]  ( .D(n2359), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[22] ) );
  DFFRHQ \uut/in2_32_reg_reg[21]  ( .D(n2358), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[21] ) );
  DFFRHQ \uut/in2_32_reg_reg[20]  ( .D(n2357), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[20] ) );
  DFFRHQ \uut/in2_32_reg_reg[19]  ( .D(n2356), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[19] ) );
  DFFRHQ \uut/in2_32_reg_reg[18]  ( .D(n2355), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[18] ) );
  DFFRHQ \uut/in2_32_reg_reg[17]  ( .D(n2354), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[17] ) );
  DFFRHQ \uut/in2_32_reg_reg[16]  ( .D(n2353), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[16] ) );
  DFFRHQ \uut/in2_32_reg_reg[15]  ( .D(n2352), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[15] ) );
  DFFRHQ \uut/in2_32_reg_reg[14]  ( .D(n2351), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[14] ) );
  DFFRHQ \uut/in2_32_reg_reg[13]  ( .D(n2350), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[13] ) );
  DFFRHQ \uut/in2_32_reg_reg[12]  ( .D(n2349), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[12] ) );
  DFFRHQ \uut/in2_32_reg_reg[11]  ( .D(n2348), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[11] ) );
  DFFRHQ \uut/in2_32_reg_reg[10]  ( .D(n2347), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[10] ) );
  DFFRHQ \uut/in2_32_reg_reg[9]  ( .D(n2346), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[9] ) );
  DFFRHQ \uut/in2_32_reg_reg[8]  ( .D(n2345), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[8] ) );
  DFFRHQ \uut/in2_32_reg_reg[7]  ( .D(n2344), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[7] ) );
  DFFRHQ \uut/in2_32_reg_reg[6]  ( .D(n2343), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[6] ) );
  DFFRHQ \uut/in2_32_reg_reg[5]  ( .D(n2342), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[5] ) );
  DFFRHQ \uut/in2_32_reg_reg[4]  ( .D(n2341), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[4] ) );
  DFFRHQ \uut/in2_32_reg_reg[3]  ( .D(n2340), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[3] ) );
  DFFRHQ \uut/in2_32_reg_reg[2]  ( .D(n2339), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[2] ) );
  DFFRHQ \uut/in2_32_reg_reg[1]  ( .D(n2338), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[1] ) );
  DFFRHQ \uut/in2_32_reg_reg[0]  ( .D(n2337), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_32_reg[0] ) );
  DFFRHQ \uut/in1_16_reg_reg[15]  ( .D(n2336), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_16_reg[15] ) );
  DFFRHQ \uut/in1_16_reg_reg[14]  ( .D(n2335), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_16_reg[14] ) );
  DFFRHQ \uut/in1_16_reg_reg[13]  ( .D(n2334), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_16_reg[13] ) );
  DFFRHQ \uut/in1_16_reg_reg[12]  ( .D(n2333), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_16_reg[12] ) );
  DFFRHQ \uut/in1_16_reg_reg[11]  ( .D(n2332), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_16_reg[11] ) );
  DFFRHQ \uut/in1_16_reg_reg[10]  ( .D(n2331), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_16_reg[10] ) );
  DFFRHQ \uut/in1_16_reg_reg[9]  ( .D(n2330), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_16_reg[9] ) );
  DFFRHQ \uut/in1_16_reg_reg[8]  ( .D(n2329), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_16_reg[8] ) );
  DFFRHQ \uut/in1_16_reg_reg[7]  ( .D(n2328), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_16_reg[7] ) );
  DFFRHQ \uut/in1_16_reg_reg[6]  ( .D(n2327), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_16_reg[6] ) );
  DFFRHQ \uut/in1_16_reg_reg[5]  ( .D(n2326), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_16_reg[5] ) );
  DFFRHQ \uut/in1_16_reg_reg[4]  ( .D(n2325), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_16_reg[4] ) );
  DFFRHQ \uut/in1_16_reg_reg[3]  ( .D(n2324), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_16_reg[3] ) );
  DFFRHQ \uut/in1_16_reg_reg[2]  ( .D(n2323), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_16_reg[2] ) );
  DFFRHQ \uut/in1_16_reg_reg[1]  ( .D(n2322), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_16_reg[1] ) );
  DFFRHQ \uut/in1_16_reg_reg[0]  ( .D(n2321), .CK(clk), .RN(rst_n), .Q(
        \uut/in1_16_reg[0] ) );
  DFFRHQ \uut/in2_16_reg_reg[15]  ( .D(n2320), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_16_reg[15] ) );
  DFFRHQ \uut/in2_16_reg_reg[14]  ( .D(n2319), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_16_reg[14] ) );
  DFFRHQ \uut/in2_16_reg_reg[13]  ( .D(n2318), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_16_reg[13] ) );
  DFFRHQ \uut/in2_16_reg_reg[12]  ( .D(n2317), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_16_reg[12] ) );
  DFFRHQ \uut/in2_16_reg_reg[11]  ( .D(n2316), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_16_reg[11] ) );
  DFFRHQ \uut/in2_16_reg_reg[10]  ( .D(n2315), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_16_reg[10] ) );
  DFFRHQ \uut/in2_16_reg_reg[9]  ( .D(n2314), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_16_reg[9] ) );
  DFFRHQ \uut/in2_16_reg_reg[8]  ( .D(n2313), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_16_reg[8] ) );
  DFFRHQ \uut/in2_16_reg_reg[7]  ( .D(n2312), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_16_reg[7] ) );
  DFFRHQ \uut/in2_16_reg_reg[6]  ( .D(n2311), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_16_reg[6] ) );
  DFFRHQ \uut/in2_16_reg_reg[5]  ( .D(n2310), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_16_reg[5] ) );
  DFFRHQ \uut/in2_16_reg_reg[4]  ( .D(n2309), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_16_reg[4] ) );
  DFFRHQ \uut/in2_16_reg_reg[3]  ( .D(n2308), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_16_reg[3] ) );
  DFFRHQ \uut/in2_16_reg_reg[2]  ( .D(n2307), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_16_reg[2] ) );
  DFFRHQ \uut/in2_16_reg_reg[1]  ( .D(n2306), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_16_reg[1] ) );
  DFFRHQ \uut/in2_16_reg_reg[0]  ( .D(n2305), .CK(clk), .RN(rst_n), .Q(
        \uut/in2_16_reg[0] ) );
  DFFRHQ \uut/start_reg  ( .D(\uut/N66 ), .CK(clk), .RN(rst_n), .Q(\uut/start ) );
  DFFRHQ \uut/mult_mant/mult8_cnt_reg[0]  ( .D(n4880), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/mult8_cnt[0] ) );
  DFFRHQ \uut/mult_mant/mult8_cnt_reg[1]  ( .D(n2484), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/mult8_cnt[1] ) );
  DFFRHQ \uut/mult_mant/mult8_cnt_reg[2]  ( .D(n2483), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/mult8_cnt[2] ) );
  DFFRHQ \uut/mult_mant/mult8_cnt_reg[3]  ( .D(n2482), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/mult8_cnt[3] ) );
  DFFRHQ \uut/mult_mant/shift_amount_reg[5]  ( .D(n2479), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/shift_amount [5]) );
  DFFRHQ \uut/mult_mant/shift_amount_reg[4]  ( .D(n2480), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/shift_amount [4]) );
  DFFRHQ \uut/mult_mant/shift_amount_reg[3]  ( .D(n2481), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/shift_amount [3]) );
  DFFRHQ \uut/mult_mant/in1_reg_reg[0]  ( .D(n4886), .CK(clk), .RN(rst_n), .Q(
        \uut/mult_mant/c1 [0]) );
  DFFRHQ \uut/mult_mant/in1_reg_reg[1]  ( .D(n4887), .CK(clk), .RN(rst_n), .Q(
        \uut/mult_mant/c1 [1]) );
  DFFRHQ \uut/mult_mant/in1_reg_reg[2]  ( .D(n4888), .CK(clk), .RN(rst_n), .Q(
        \uut/mult_mant/c1 [2]) );
  DFFRHQ \uut/mult_mant/in1_reg_reg[3]  ( .D(n4889), .CK(clk), .RN(rst_n), .Q(
        \uut/mult_mant/c1 [3]) );
  DFFRHQ \uut/mult_mant/in1_reg_reg[4]  ( .D(n4890), .CK(clk), .RN(rst_n), .Q(
        \uut/mult_mant/c1 [4]) );
  DFFRHQ \uut/mult_mant/in1_reg_reg[5]  ( .D(n4891), .CK(clk), .RN(rst_n), .Q(
        \uut/mult_mant/c1 [5]) );
  DFFRHQ \uut/mult_mant/in1_reg_reg[6]  ( .D(n4892), .CK(clk), .RN(rst_n), .Q(
        \uut/mult_mant/c1 [6]) );
  DFFRHQ \uut/mult_mant/in1_reg_reg[7]  ( .D(n4893), .CK(clk), .RN(rst_n), .Q(
        \uut/mult_mant/c1 [7]) );
  DFFRHQ \uut/mult_mant/in1_reg_reg[8]  ( .D(n4894), .CK(clk), .RN(rst_n), .Q(
        \uut/mult_mant/b1 [0]) );
  DFFRHQ \uut/mult_mant/in1_reg_reg[9]  ( .D(n4895), .CK(clk), .RN(rst_n), .Q(
        \uut/mult_mant/b1 [1]) );
  DFFRHQ \uut/mult_mant/in1_reg_reg[10]  ( .D(n4896), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/b1 [2]) );
  DFFRHQ \uut/mult_mant/in1_reg_reg[11]  ( .D(n2293), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/b1 [3]) );
  DFFRHQ \uut/mult_mant/in1_reg_reg[12]  ( .D(n2292), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/b1 [4]) );
  DFFRHQ \uut/mult_mant/in1_reg_reg[13]  ( .D(n2291), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/b1 [5]) );
  DFFRHQ \uut/mult_mant/in1_reg_reg[14]  ( .D(n2290), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/b1 [6]) );
  DFFRHQ \uut/mult_mant/in1_reg_reg[15]  ( .D(n2289), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/b1 [7]) );
  DFFRHQ \uut/mult_mant/in1_reg_reg[16]  ( .D(n2288), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/a1 [0]) );
  DFFRHQ \uut/mult_mant/in1_segment_reg[0]  ( .D(n2478), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/in1_segment [0]) );
  DFFRHQ \uut/mult_mant/in1_reg_reg[17]  ( .D(n2287), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/a1 [1]) );
  DFFRHQ \uut/mult_mant/in1_segment_reg[1]  ( .D(n2477), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/in1_segment [1]) );
  DFFRHQ \uut/mult_mant/in1_reg_reg[18]  ( .D(n2286), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/a1 [2]) );
  DFFRHQ \uut/mult_mant/in1_segment_reg[2]  ( .D(n2476), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/in1_segment [2]) );
  DFFRHQ \uut/mult_mant/in1_reg_reg[19]  ( .D(n2285), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/a1 [3]) );
  DFFRHQ \uut/mult_mant/in1_segment_reg[3]  ( .D(n2475), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/in1_segment [3]) );
  DFFRHQ \uut/mult_mant/in1_reg_reg[20]  ( .D(n2284), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/a1 [4]) );
  DFFRHQ \uut/mult_mant/in1_segment_reg[4]  ( .D(n2474), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/in1_segment [4]) );
  DFFRHQ \uut/mult_mant/in1_reg_reg[21]  ( .D(n2283), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/a1 [5]) );
  DFFRHQ \uut/mult_mant/in1_segment_reg[5]  ( .D(n2473), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/in1_segment [5]) );
  DFFRHQ \uut/mult_mant/in1_reg_reg[22]  ( .D(n2282), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/a1 [6]) );
  DFFRHQ \uut/mult_mant/in1_segment_reg[6]  ( .D(n2472), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/in1_segment [6]) );
  DFFRHQ \uut/mult_mant/in1_reg_reg[23]  ( .D(n2281), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/a1 [7]) );
  DFFRHQ \uut/mult_mant/in1_segment_reg[7]  ( .D(n2471), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/in1_segment [7]) );
  DFFRHQ \uut/mult_mant/in2_reg_reg[0]  ( .D(n4897), .CK(clk), .RN(rst_n), .Q(
        \uut/mult_mant/c2 [0]) );
  DFFRHQ \uut/mult_mant/in2_reg_reg[1]  ( .D(n4898), .CK(clk), .RN(rst_n), .Q(
        \uut/mult_mant/c2 [1]) );
  DFFRHQ \uut/mult_mant/in2_reg_reg[2]  ( .D(n4899), .CK(clk), .RN(rst_n), .Q(
        \uut/mult_mant/c2 [2]) );
  DFFRHQ \uut/mult_mant/in2_reg_reg[3]  ( .D(n4900), .CK(clk), .RN(rst_n), .Q(
        \uut/mult_mant/c2 [3]) );
  DFFRHQ \uut/mult_mant/in2_reg_reg[4]  ( .D(n4901), .CK(clk), .RN(rst_n), .Q(
        \uut/mult_mant/c2 [4]) );
  DFFRHQ \uut/mult_mant/in2_reg_reg[5]  ( .D(n4902), .CK(clk), .RN(rst_n), .Q(
        \uut/mult_mant/c2 [5]) );
  DFFRHQ \uut/mult_mant/in2_reg_reg[6]  ( .D(n4903), .CK(clk), .RN(rst_n), .Q(
        \uut/mult_mant/c2 [6]) );
  DFFRHQ \uut/mult_mant/in2_reg_reg[7]  ( .D(n4904), .CK(clk), .RN(rst_n), .Q(
        \uut/mult_mant/c2 [7]) );
  DFFRHQ \uut/mult_mant/in2_reg_reg[8]  ( .D(n4905), .CK(clk), .RN(rst_n), .Q(
        \uut/mult_mant/b2 [0]) );
  DFFRHQ \uut/mult_mant/in2_reg_reg[9]  ( .D(n4906), .CK(clk), .RN(rst_n), .Q(
        \uut/mult_mant/b2 [1]) );
  DFFRHQ \uut/mult_mant/in2_reg_reg[10]  ( .D(n4907), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/b2 [2]) );
  DFFRHQ \uut/mult_mant/in2_reg_reg[11]  ( .D(n2269), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/b2 [3]) );
  DFFRHQ \uut/mult_mant/in2_reg_reg[12]  ( .D(n2268), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/b2 [4]) );
  DFFRHQ \uut/mult_mant/in2_reg_reg[13]  ( .D(n2267), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/b2 [5]) );
  DFFRHQ \uut/mult_mant/in2_reg_reg[14]  ( .D(n2266), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/b2 [6]) );
  DFFRHQ \uut/mult_mant/in2_reg_reg[15]  ( .D(n2265), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/b2 [7]) );
  DFFRHQ \uut/mult_mant/in2_reg_reg[16]  ( .D(n2264), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/a2 [0]) );
  DFFRHQ \uut/mult_mant/in2_segment_reg[0]  ( .D(n2470), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/in2_segment [0]) );
  DFFRHQ \uut/mult_mant/in2_reg_reg[17]  ( .D(n2263), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/a2 [1]) );
  DFFRHQ \uut/mult_mant/in2_segment_reg[1]  ( .D(n2469), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/in2_segment [1]) );
  DFFRHQ \uut/mult_mant/in2_reg_reg[18]  ( .D(n2262), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/a2 [2]) );
  DFFRHQ \uut/mult_mant/in2_segment_reg[2]  ( .D(n2468), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/in2_segment [2]) );
  DFFRHQ \uut/mult_mant/in2_reg_reg[19]  ( .D(n2261), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/a2 [3]) );
  DFFRHQ \uut/mult_mant/in2_segment_reg[3]  ( .D(n2467), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/in2_segment [3]) );
  DFFRHQ \uut/mult_mant/in2_reg_reg[20]  ( .D(n2260), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/a2 [4]) );
  DFFRHQ \uut/mult_mant/in2_segment_reg[4]  ( .D(n2466), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/in2_segment [4]) );
  DFFRHQ \uut/mult_mant/in2_reg_reg[21]  ( .D(n2259), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/a2 [5]) );
  DFFRHQ \uut/mult_mant/in2_segment_reg[5]  ( .D(n2465), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/in2_segment [5]) );
  DFFRHQ \uut/mult_mant/in2_reg_reg[22]  ( .D(n2258), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/a2 [6]) );
  DFFRHQ \uut/mult_mant/in2_segment_reg[6]  ( .D(n2464), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/in2_segment [6]) );
  DFFRHQ \uut/mult_mant/in2_reg_reg[23]  ( .D(n2257), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/a2 [7]) );
  DFFRHQ \uut/mult_mant/in2_segment_reg[7]  ( .D(n2463), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/in2_segment [7]) );
  DFFRHQ \uut/mult_mant/temp_product_reg[47]  ( .D(n4960), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[47] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[46]  ( .D(n4959), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[46] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[45]  ( .D(n4913), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[45] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[44]  ( .D(n4914), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[44] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[43]  ( .D(n4915), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[43] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[42]  ( .D(n4916), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[42] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[41]  ( .D(n4917), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[41] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[40]  ( .D(n4918), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[40] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[39]  ( .D(n4919), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[39] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[38]  ( .D(n4920), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[38] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[37]  ( .D(n4921), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[37] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[36]  ( .D(n4922), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[36] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[35]  ( .D(n4923), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[35] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[34]  ( .D(n4924), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[34] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[33]  ( .D(n4925), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[33] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[32]  ( .D(n4926), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[32] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[31]  ( .D(n4927), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[31] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[30]  ( .D(n4928), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[30] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[29]  ( .D(n4929), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[29] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[28]  ( .D(n4930), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[28] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[27]  ( .D(n4931), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[27] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[26]  ( .D(n4932), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[26] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[25]  ( .D(n4933), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[25] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[24]  ( .D(n4934), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[24] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[23]  ( .D(n4935), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[23] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[22]  ( .D(n4936), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[22] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[21]  ( .D(n4937), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[21] ) );
  DFFRHQ \uut/mult_mant/normalize_reg  ( .D(n2462), .CK(clk), .RN(rst_n), .Q(
        \uut/normalize ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[20]  ( .D(n4938), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[20] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[19]  ( .D(n4939), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[19] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[18]  ( .D(n4940), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[18] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[17]  ( .D(n4941), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[17] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[16]  ( .D(n4942), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[16] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[15]  ( .D(n4943), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[15] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[14]  ( .D(n4944), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[14] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[13]  ( .D(n4945), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[13] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[12]  ( .D(n4946), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[12] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[11]  ( .D(n4947), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[11] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[10]  ( .D(n4948), .CK(clk), .RN(rst_n), .Q(\uut/mult_mant/temp_product[10] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[9]  ( .D(n4949), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/temp_product[9] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[8]  ( .D(n4950), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/temp_product[8] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[7]  ( .D(n4951), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/temp_product[7] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[6]  ( .D(n4952), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/temp_product[6] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[5]  ( .D(n4953), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/temp_product[5] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[4]  ( .D(n4954), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/temp_product[4] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[3]  ( .D(n4955), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/temp_product[3] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[2]  ( .D(n4956), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/temp_product[2] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[1]  ( .D(n4957), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/temp_product[1] ) );
  DFFRHQ \uut/mult_mant/temp_product_reg[0]  ( .D(n4958), .CK(clk), .RN(rst_n), 
        .Q(\uut/mult_mant/temp_product[0] ) );
  DFFRHQ \uut/mult_mant/product_reg[0]  ( .D(n2256), .CK(clk), .RN(rst_n), .Q(
        \uut/mant_out[0] ) );
  DFFRHQ \uut/mult_mant/product_reg[1]  ( .D(n2255), .CK(clk), .RN(rst_n), .Q(
        \uut/mant_out[1] ) );
  DFFRHQ \uut/mult_mant/product_reg[2]  ( .D(n2254), .CK(clk), .RN(rst_n), .Q(
        \uut/mant_out[2] ) );
  DFFRHQ \uut/mult_mant/product_reg[3]  ( .D(n2253), .CK(clk), .RN(rst_n), .Q(
        \uut/mant_out[3] ) );
  DFFRHQ \bit0_reg[0]  ( .D(N5258), .CK(clk), .RN(rst_n), .Q(bit0[0]) );
  DFFRHQ \bit0_reg[1]  ( .D(N5259), .CK(clk), .RN(rst_n), .Q(bit0[1]) );
  DFFRHQ \bit0_reg[4]  ( .D(N5262), .CK(clk), .RN(rst_n), .Q(bit0[4]) );
  DFFRHQ \bit0_reg[2]  ( .D(N5260), .CK(clk), .RN(rst_n), .Q(bit0[2]) );
  DFFRHQ \bit0_reg[6]  ( .D(N5264), .CK(clk), .RN(rst_n), .Q(bit0[6]) );
  DFFRHQ \bit0_reg[5]  ( .D(N5263), .CK(clk), .RN(rst_n), .Q(bit0[5]) );
  DFFRHQ \bit0_reg[3]  ( .D(N5261), .CK(clk), .RN(rst_n), .Q(bit0[3]) );
  DFFRHQ \uut/mult_mant/product_reg[4]  ( .D(n2252), .CK(clk), .RN(rst_n), .Q(
        \uut/mant_out[4] ) );
  DFFRHQ \uut/mult_mant/product_reg[5]  ( .D(n2251), .CK(clk), .RN(rst_n), .Q(
        \uut/mant_out[5] ) );
  DFFRHQ \uut/mult_mant/product_reg[6]  ( .D(n2250), .CK(clk), .RN(rst_n), .Q(
        \uut/mant_out[6] ) );
  DFFRHQ \uut/mult_mant/product_reg[7]  ( .D(n2249), .CK(clk), .RN(rst_n), .Q(
        \uut/mant_out[7] ) );
  DFFRHQ \bit1_reg[0]  ( .D(N5144), .CK(clk), .RN(rst_n), .Q(bit1[0]) );
  DFFRHQ \bit1_reg[1]  ( .D(N5145), .CK(clk), .RN(rst_n), .Q(bit1[1]) );
  DFFRHQ \bit1_reg[4]  ( .D(N5148), .CK(clk), .RN(rst_n), .Q(bit1[4]) );
  DFFRHQ \bit1_reg[2]  ( .D(N5146), .CK(clk), .RN(rst_n), .Q(bit1[2]) );
  DFFRHQ \bit1_reg[6]  ( .D(N5150), .CK(clk), .RN(rst_n), .Q(bit1[6]) );
  DFFRHQ \bit1_reg[5]  ( .D(N5149), .CK(clk), .RN(rst_n), .Q(bit1[5]) );
  DFFRHQ \bit1_reg[3]  ( .D(N5147), .CK(clk), .RN(rst_n), .Q(bit1[3]) );
  DFFRHQ \uut/mult_mant/product_reg[8]  ( .D(n2248), .CK(clk), .RN(rst_n), .Q(
        \uut/mant_out[8] ) );
  DFFRHQ \uut/mult_mant/product_reg[9]  ( .D(n2247), .CK(clk), .RN(rst_n), .Q(
        \uut/mant_out[9] ) );
  DFFRHQ \uut/mult_mant/product_reg[10]  ( .D(n2246), .CK(clk), .RN(rst_n), 
        .Q(\uut/mant_out[10] ) );
  DFFRHQ \uut/mult_mant/product_reg[11]  ( .D(n2245), .CK(clk), .RN(rst_n), 
        .Q(\uut/mant_out[11] ) );
  DFFRHQ \uut/mult_mant/product_reg[12]  ( .D(n2244), .CK(clk), .RN(rst_n), 
        .Q(\uut/mant_out[12] ) );
  DFFRHQ \uut/mult_mant/product_reg[13]  ( .D(n2243), .CK(clk), .RN(rst_n), 
        .Q(\uut/mant_out[13] ) );
  DFFRHQ \uut/mult_mant/product_reg[14]  ( .D(n2242), .CK(clk), .RN(rst_n), 
        .Q(\uut/mant_out[14] ) );
  DFFRHQ \uut/mult_mant/product_reg[15]  ( .D(n2241), .CK(clk), .RN(rst_n), 
        .Q(\uut/mant_out[15] ) );
  DFFRHQ \uut/mult_mant/product_reg[16]  ( .D(n2240), .CK(clk), .RN(rst_n), 
        .Q(\uut/mant_out[16] ) );
  DFFRHQ \uut/mult_mant/product_reg[17]  ( .D(n2239), .CK(clk), .RN(rst_n), 
        .Q(\uut/mant_out[17] ) );
  DFFRHQ \uut/mult_mant/product_reg[18]  ( .D(n2238), .CK(clk), .RN(rst_n), 
        .Q(\uut/mant_out[18] ) );
  DFFRHQ \uut/mult_mant/product_reg[19]  ( .D(n2237), .CK(clk), .RN(rst_n), 
        .Q(\uut/mant_out[19] ) );
  DFFRHQ \bit4_reg[2]  ( .D(N4804), .CK(clk), .RN(rst_n), .Q(bit4[2]) );
  DFFRHQ \bit4_reg[1]  ( .D(N4803), .CK(clk), .RN(rst_n), .Q(bit4[1]) );
  DFFRHQ \bit4_reg[4]  ( .D(N4806), .CK(clk), .RN(rst_n), .Q(bit4[4]) );
  DFFRHQ \bit4_reg[5]  ( .D(N4807), .CK(clk), .RN(rst_n), .Q(bit4[5]) );
  DFFRHQ \bit4_reg[0]  ( .D(N4802), .CK(clk), .RN(rst_n), .Q(bit4[0]) );
  DFFRHQ \bit4_reg[6]  ( .D(N4808), .CK(clk), .RN(rst_n), .Q(bit4[6]) );
  DFFRHQ \bit4_reg[3]  ( .D(N4805), .CK(clk), .RN(rst_n), .Q(bit4[3]) );
  DFFRHQ \uut/mult_mant/product_reg[20]  ( .D(n2236), .CK(clk), .RN(rst_n), 
        .Q(\uut/mant_out[20] ) );
  DFFRHQ \uut/mult_mant/product_reg[21]  ( .D(n2235), .CK(clk), .RN(rst_n), 
        .Q(\uut/mant_out[21] ) );
  DFFRHQ \uut/mult_mant/product_reg[22]  ( .D(n2234), .CK(clk), .RN(rst_n), 
        .Q(\uut/mant_out[22] ) );
  DFFRHQ \uut/mult_mant/more_than_1_reg  ( .D(n2461), .CK(clk), .RN(rst_n), 
        .Q(\uut/more_than_1 ) );
  DFFRHQ \uut/exp_complete_reg  ( .D(n4912), .CK(clk), .RN(rst_n), .Q(
        \uut/exp_complete ) );
  DFFRHQ \uut/exp_out_reg[8]  ( .D(n4881), .CK(clk), .RN(rst_n), .Q(
        \uut/exp_out[8] ) );
  DFFRHQ \uut/exp_out_reg[7]  ( .D(n4882), .CK(clk), .RN(rst_n), .Q(
        \uut/exp_out[7] ) );
  DFFRHQ \uut/exp_out_reg[6]  ( .D(n4883), .CK(clk), .RN(rst_n), .Q(
        \uut/exp_out[6] ) );
  DFFRHQ \uut/exp_out_reg[5]  ( .D(n4884), .CK(clk), .RN(rst_n), .Q(
        \uut/exp_out[5] ) );
  DFFRHQ \bit7_reg[6]  ( .D(N4622), .CK(clk), .RN(rst_n), .Q(bit7[6]) );
  DFFRHQ \bit7_reg[2]  ( .D(N4618), .CK(clk), .RN(rst_n), .Q(bit7[2]) );
  DFFRHQ \bit7_reg[1]  ( .D(N4617), .CK(clk), .RN(rst_n), .Q(bit7[1]) );
  DFFRHQ \bit7_reg[0]  ( .D(N4616), .CK(clk), .RN(rst_n), .Q(bit7[0]) );
  DFFRHQ \bit7_reg[5]  ( .D(N4621), .CK(clk), .RN(rst_n), .Q(bit7[5]) );
  DFFRHQ \bit7_reg[4]  ( .D(N4620), .CK(clk), .RN(rst_n), .Q(bit7[4]) );
  DFFRHQ \bit7_reg[3]  ( .D(N4619), .CK(clk), .RN(rst_n), .Q(bit7[3]) );
  DFFRHQ \uut/exp_out_reg[4]  ( .D(n4885), .CK(clk), .RN(rst_n), .Q(
        \uut/exp_out[4] ) );
  DFFRHQ \uut/exp_out_reg[3]  ( .D(n4909), .CK(clk), .RN(rst_n), .Q(
        \uut/exp_out[3] ) );
  DFFRHQ \uut/exp_out_reg[2]  ( .D(n4910), .CK(clk), .RN(rst_n), .Q(
        \uut/exp_out[2] ) );
  DFFRHQ \bit3_reg[0]  ( .D(N4916), .CK(clk), .RN(rst_n), .Q(bit3[0]) );
  DFFRHQ \bit3_reg[3]  ( .D(N4919), .CK(clk), .RN(rst_n), .Q(bit3[3]) );
  DFFRHQ \bit3_reg[4]  ( .D(N4920), .CK(clk), .RN(rst_n), .Q(bit3[4]) );
  DFFRHQ \bit3_reg[6]  ( .D(N4922), .CK(clk), .RN(rst_n), .Q(bit3[6]) );
  DFFRHQ \bit3_reg[5]  ( .D(N4921), .CK(clk), .RN(rst_n), .Q(bit3[5]) );
  DFFRHQ \bit3_reg[2]  ( .D(N4918), .CK(clk), .RN(rst_n), .Q(bit3[2]) );
  DFFRHQ \bit3_reg[1]  ( .D(N4917), .CK(clk), .RN(rst_n), .Q(bit3[1]) );
  DFFRHQ \uut/exp_out_reg[1]  ( .D(n4911), .CK(clk), .RN(rst_n), .Q(
        \uut/exp_out[1] ) );
  DFFRHQ \bit6_reg[6]  ( .D(N4684), .CK(clk), .RN(rst_n), .Q(bit6[6]) );
  DFFRHQ \bit6_reg[2]  ( .D(N4680), .CK(clk), .RN(rst_n), .Q(bit6[2]) );
  DFFRHQ \bit6_reg[1]  ( .D(N4679), .CK(clk), .RN(rst_n), .Q(bit6[1]) );
  DFFRHQ \bit6_reg[0]  ( .D(N4678), .CK(clk), .RN(rst_n), .Q(bit6[0]) );
  DFFRHQ \bit6_reg[4]  ( .D(N4682), .CK(clk), .RN(rst_n), .Q(bit6[4]) );
  DFFRHQ \bit6_reg[5]  ( .D(N4683), .CK(clk), .RN(rst_n), .Q(bit6[5]) );
  DFFRHQ \bit6_reg[3]  ( .D(N4681), .CK(clk), .RN(rst_n), .Q(bit6[3]) );
  DFFRHQ \uut/exp_out_reg[0]  ( .D(n4908), .CK(clk), .RN(rst_n), .Q(
        \uut/exp_out[0] ) );
  DFFRHQ \bit5_reg[2]  ( .D(N4742), .CK(clk), .RN(rst_n), .Q(bit5[2]) );
  DFFRHQ \bit5_reg[1]  ( .D(N4741), .CK(clk), .RN(rst_n), .Q(bit5[1]) );
  DFFRHQ \bit5_reg[4]  ( .D(N4744), .CK(clk), .RN(rst_n), .Q(bit5[4]) );
  DFFRHQ \bit5_reg[5]  ( .D(N4745), .CK(clk), .RN(rst_n), .Q(bit5[5]) );
  DFFRHQ \bit5_reg[0]  ( .D(N4740), .CK(clk), .RN(rst_n), .Q(bit5[0]) );
  DFFRHQ \bit5_reg[6]  ( .D(N4746), .CK(clk), .RN(rst_n), .Q(bit5[6]) );
  DFFRHQ \bit5_reg[3]  ( .D(N4743), .CK(clk), .RN(rst_n), .Q(bit5[3]) );
  DFFRHQ \bit2_reg[2]  ( .D(N5032), .CK(clk), .RN(rst_n), .Q(bit2[2]) );
  DFFRHQ \bit2_reg[4]  ( .D(N5034), .CK(clk), .RN(rst_n), .Q(bit2[4]) );
  DFFRHQ \bit2_reg[3]  ( .D(N5033), .CK(clk), .RN(rst_n), .Q(bit2[3]) );
  DFFRHQ \bit2_reg[5]  ( .D(N5035), .CK(clk), .RN(rst_n), .Q(bit2[5]) );
  DFFRHQ \bit2_reg[6]  ( .D(N5036), .CK(clk), .RN(rst_n), .Q(bit2[6]) );
  DFFRHQ \bit2_reg[0]  ( .D(N5030), .CK(clk), .RN(rst_n), .Q(bit2[0]) );
  DFFRHQ \bit2_reg[1]  ( .D(N5031), .CK(clk), .RN(rst_n), .Q(bit2[1]) );
  OR2 U2826 ( .A(n2769), .B(ce), .Y(n2518) );
  OR2 U2827 ( .A(n2771), .B(ce), .Y(n2519) );
  OR2 U2828 ( .A(data_type), .B(n2788), .Y(n2520) );
  OR3 U2829 ( .A(\uut/mult_mant/mult8_cnt[1] ), .B(
        \uut/mult_mant/mult8_cnt[3] ), .C(n3520), .Y(n2521) );
  OR2 U2830 ( .A(error), .B(n2734), .Y(n2522) );
  OR2 U2831 ( .A(n3755), .B(n2734), .Y(n2523) );
  OR2 U2832 ( .A(n3827), .B(n2734), .Y(n2524) );
  OR3 U2833 ( .A(\uut/mult_mant/mult8_cnt[3] ), .B(n3520), .C(n3452), .Y(n2525) );
  OR2 U2834 ( .A(n4773), .B(n2770), .Y(n2526) );
  OR2 U2835 ( .A(n4858), .B(n2772), .Y(n2527) );
  AND2 U2836 ( .A(n3391), .B(\uut/mult_mant/state[1] ), .Y(n2528) );
  AND2 U2837 ( .A(ready), .B(enter), .Y(n2529) );
  AND2 U2838 ( .A(\uut/start ), .B(data_type), .Y(n2530) );
  NOR2 U2839 ( .A(data_type), .B(enter), .Y(n2531) );
  INV U2840 ( .A(n2858), .Y(n2532) );
  INV U2841 ( .A(n2532), .Y(n2533) );
  INV U2842 ( .A(n4095), .Y(n2534) );
  INV U2843 ( .A(n2534), .Y(n2535) );
  INV U2844 ( .A(n3594), .Y(n2536) );
  INV U2845 ( .A(n2536), .Y(n2537) );
  INV U2846 ( .A(\uut/exp_complete ), .Y(n2538) );
  INV U2847 ( .A(n2538), .Y(n2539) );
  INV U2848 ( .A(\uut/mult_mant/mult8_cnt[0] ), .Y(n2540) );
  INV U2849 ( .A(n2540), .Y(n2541) );
  INV U2850 ( .A(n4016), .Y(n2542) );
  INV U2851 ( .A(n2542), .Y(n2543) );
  INV U2852 ( .A(n2530), .Y(n2544) );
  INV U2853 ( .A(n2530), .Y(n2545) );
  INV U2854 ( .A(n3895), .Y(n2546) );
  INV U2855 ( .A(n2546), .Y(n2547) );
  INV U2856 ( .A(\uut/mult_mant/shift_amount [4]), .Y(n2548) );
  INV U2857 ( .A(n2548), .Y(n2549) );
  INV U2858 ( .A(n3913), .Y(n2550) );
  INV U2859 ( .A(n2550), .Y(n2551) );
  INV U2860 ( .A(n3917), .Y(n2552) );
  INV U2861 ( .A(n2552), .Y(n2553) );
  INV U2862 ( .A(n3977), .Y(n2554) );
  INV U2863 ( .A(n2554), .Y(n2555) );
  INV U2864 ( .A(n4036), .Y(n2556) );
  INV U2865 ( .A(n2556), .Y(n2557) );
  INV U2866 ( .A(n3449), .Y(n2558) );
  INV U2867 ( .A(n2558), .Y(n2559) );
  INV U2868 ( .A(n3439), .Y(n2560) );
  INV U2869 ( .A(n2560), .Y(n2561) );
  INV U2870 ( .A(n5002), .Y(n2562) );
  INV U2871 ( .A(n2562), .Y(out_sel[5]) );
  INV U2872 ( .A(n5004), .Y(n2564) );
  INV U2873 ( .A(n2564), .Y(out_sel[3]) );
  INV U2874 ( .A(n5003), .Y(n2566) );
  INV U2875 ( .A(n2566), .Y(out_sel[4]) );
  INV U2876 ( .A(n5006), .Y(n2568) );
  INV U2877 ( .A(n2568), .Y(out_sel[1]) );
  INV U2878 ( .A(n5005), .Y(n2570) );
  INV U2879 ( .A(n2570), .Y(out_sel[2]) );
  INV U2880 ( .A(n4996), .Y(n2572) );
  INV U2881 ( .A(n2572), .Y(disp2_sel[5]) );
  INV U2882 ( .A(n4995), .Y(n2574) );
  INV U2883 ( .A(n2574), .Y(disp2_sel[6]) );
  INV U2884 ( .A(n4997), .Y(n2576) );
  INV U2885 ( .A(n2576), .Y(disp2_sel[4]) );
  INV U2886 ( .A(n5000), .Y(n2578) );
  INV U2887 ( .A(n2578), .Y(disp2_sel[1]) );
  INV U2888 ( .A(n4999), .Y(n2580) );
  INV U2889 ( .A(n2580), .Y(disp2_sel[2]) );
  INV U2890 ( .A(n4990), .Y(n2582) );
  INV U2891 ( .A(n2582), .Y(disp1_sel[5]) );
  INV U2892 ( .A(n4989), .Y(n2584) );
  INV U2893 ( .A(n2584), .Y(disp1_sel[6]) );
  INV U2894 ( .A(n4991), .Y(n2586) );
  INV U2895 ( .A(n2586), .Y(disp1_sel[4]) );
  INV U2896 ( .A(n4994), .Y(n2588) );
  INV U2897 ( .A(n2588), .Y(disp1_sel[1]) );
  INV U2898 ( .A(n4993), .Y(n2590) );
  INV U2899 ( .A(n2590), .Y(disp1_sel[2]) );
  INV U2900 ( .A(N5398), .Y(n2592) );
  INV U2901 ( .A(n2592), .Y(out_sel[0]) );
  INV U2902 ( .A(N5346), .Y(n2594) );
  INV U2903 ( .A(n2594), .Y(disp2_sel[0]) );
  INV U2904 ( .A(N5294), .Y(n2596) );
  INV U2905 ( .A(n2596), .Y(disp1_sel[0]) );
  INV U2906 ( .A(in2_disp[31]), .Y(n2598) );
  INV U2907 ( .A(n2598), .Y(n2599) );
  INV U2908 ( .A(in2_disp[27]), .Y(n2600) );
  INV U2909 ( .A(n2600), .Y(n2601) );
  INV U2910 ( .A(in2_disp[23]), .Y(n2602) );
  INV U2911 ( .A(n2602), .Y(n2603) );
  INV U2912 ( .A(in2_disp[19]), .Y(n2604) );
  INV U2913 ( .A(n2604), .Y(n2605) );
  INV U2914 ( .A(in2_disp[12]), .Y(n2606) );
  INV U2915 ( .A(n2606), .Y(n2607) );
  INV U2916 ( .A(in2_disp[14]), .Y(n2608) );
  INV U2917 ( .A(n2608), .Y(n2609) );
  INV U2918 ( .A(in2_disp[4]), .Y(n2610) );
  INV U2919 ( .A(n2610), .Y(n2611) );
  INV U2920 ( .A(in2_disp[6]), .Y(n2612) );
  INV U2921 ( .A(n2612), .Y(n2613) );
  INV U2922 ( .A(in2_disp[0]), .Y(n2614) );
  INV U2923 ( .A(n2614), .Y(n2615) );
  INV U2924 ( .A(in2_disp[2]), .Y(n2616) );
  INV U2925 ( .A(n2616), .Y(n2617) );
  INV U2926 ( .A(in1_disp[31]), .Y(n2618) );
  INV U2927 ( .A(n2618), .Y(n2619) );
  INV U2928 ( .A(in1_disp[27]), .Y(n2620) );
  INV U2929 ( .A(n2620), .Y(n2621) );
  INV U2930 ( .A(in1_disp[23]), .Y(n2622) );
  INV U2931 ( .A(n2622), .Y(n2623) );
  INV U2932 ( .A(in1_disp[19]), .Y(n2624) );
  INV U2933 ( .A(n2624), .Y(n2625) );
  INV U2934 ( .A(in1_disp[12]), .Y(n2626) );
  INV U2935 ( .A(n2626), .Y(n2627) );
  INV U2936 ( .A(in1_disp[14]), .Y(n2628) );
  INV U2937 ( .A(n2628), .Y(n2629) );
  INV U2938 ( .A(in1_disp[4]), .Y(n2630) );
  INV U2939 ( .A(n2630), .Y(n2631) );
  INV U2940 ( .A(in1_disp[6]), .Y(n2632) );
  INV U2941 ( .A(n2632), .Y(n2633) );
  INV U2942 ( .A(in1_disp[0]), .Y(n2634) );
  INV U2943 ( .A(n2634), .Y(n2635) );
  INV U2944 ( .A(in1_disp[2]), .Y(n2636) );
  INV U2945 ( .A(n2636), .Y(n2637) );
  INV U2946 ( .A(n3847), .Y(n2638) );
  INV U2947 ( .A(n2638), .Y(n2639) );
  INV U2948 ( .A(n4988), .Y(n2640) );
  INV U2949 ( .A(n2640), .Y(n2641) );
  INV U2950 ( .A(n3190), .Y(n2642) );
  INV U2951 ( .A(n2642), .Y(n2643) );
  INV U2952 ( .A(n3206), .Y(n2644) );
  INV U2953 ( .A(n2644), .Y(n2645) );
  INV U2954 ( .A(n3694), .Y(n2646) );
  INV U2955 ( .A(n2646), .Y(n2647) );
  INV U2956 ( .A(n3766), .Y(n2648) );
  INV U2957 ( .A(n2648), .Y(n2649) );
  INV U2958 ( .A(n2526), .Y(n2650) );
  INV U2959 ( .A(n2527), .Y(n2651) );
  INV U2960 ( .A(n3475), .Y(n2652) );
  INV U2961 ( .A(n2652), .Y(n2653) );
  INV U2962 ( .A(n3474), .Y(n2654) );
  INV U2963 ( .A(n2654), .Y(n2655) );
  INV U2964 ( .A(n4714), .Y(n2656) );
  INV U2965 ( .A(n2656), .Y(n2657) );
  INV U2966 ( .A(n4799), .Y(n2658) );
  INV U2967 ( .A(n2658), .Y(n2659) );
  INV U2968 ( .A(n3476), .Y(n2660) );
  INV U2969 ( .A(n2660), .Y(n2661) );
  INV U2970 ( .A(n3496), .Y(n2662) );
  INV U2971 ( .A(n2662), .Y(n2663) );
  INV U2972 ( .A(n3907), .Y(n2664) );
  INV U2973 ( .A(n2664), .Y(n2665) );
  INV U2974 ( .A(n3969), .Y(n2666) );
  INV U2975 ( .A(n2666), .Y(n2667) );
  INV U2976 ( .A(n3999), .Y(n2668) );
  INV U2977 ( .A(n2668), .Y(n2669) );
  INV U2978 ( .A(n4028), .Y(n2670) );
  INV U2979 ( .A(n2670), .Y(n2671) );
  INV U2980 ( .A(in1_disp[20]), .Y(n2672) );
  INV U2981 ( .A(n2672), .Y(n2673) );
  INV U2982 ( .A(in1_disp[16]), .Y(n2674) );
  INV U2983 ( .A(n2674), .Y(n2675) );
  INV U2984 ( .A(in2_disp[16]), .Y(n2676) );
  INV U2985 ( .A(n2676), .Y(n2677) );
  INV U2986 ( .A(in1_disp[28]), .Y(n2678) );
  INV U2987 ( .A(n2678), .Y(n2679) );
  INV U2988 ( .A(in2_disp[28]), .Y(n2680) );
  INV U2989 ( .A(n2680), .Y(n2681) );
  INV U2990 ( .A(in2_disp[20]), .Y(n2682) );
  INV U2991 ( .A(n2682), .Y(n2683) );
  INV U2992 ( .A(n2523), .Y(n2684) );
  INV U2993 ( .A(n2524), .Y(n2685) );
  INV U2994 ( .A(n3906), .Y(n2686) );
  INV U2995 ( .A(n2686), .Y(n2687) );
  INV U2996 ( .A(n3912), .Y(n2688) );
  INV U2997 ( .A(n2688), .Y(n2689) );
  INV U2998 ( .A(n3696), .Y(n2690) );
  INV U2999 ( .A(n2690), .Y(n2691) );
  INV U3000 ( .A(n3768), .Y(n2692) );
  INV U3001 ( .A(n2692), .Y(n2693) );
  INV U3002 ( .A(n3833), .Y(n2694) );
  INV U3003 ( .A(n2694), .Y(n2695) );
  INV U3004 ( .A(n2785), .Y(n2696) );
  INV U3005 ( .A(n2696), .Y(n2697) );
  INV U3006 ( .A(\uut/mult_mant/shift_amount [3]), .Y(n2698) );
  INV U3007 ( .A(n2698), .Y(n2699) );
  INV U3008 ( .A(n3841), .Y(n2700) );
  INV U3009 ( .A(n2700), .Y(n2701) );
  INV U3010 ( .A(N5271), .Y(n2702) );
  INV U3011 ( .A(n2702), .Y(disp1_sel[7]) );
  INV U3012 ( .A(n2522), .Y(n2704) );
  INV U3013 ( .A(n4987), .Y(n2705) );
  INV U3014 ( .A(n2705), .Y(out_sel[7]) );
  INV U3015 ( .A(N5323), .Y(n2707) );
  INV U3016 ( .A(n2707), .Y(disp2_sel[7]) );
  INV U3017 ( .A(n4064), .Y(n2709) );
  INV U3018 ( .A(n2709), .Y(n2710) );
  INV U3019 ( .A(n5001), .Y(n2711) );
  INV U3020 ( .A(n2711), .Y(out_sel[6]) );
  INV U3021 ( .A(n2525), .Y(n2713) );
  INV U3022 ( .A(n3836), .Y(n2714) );
  INV U3023 ( .A(n2714), .Y(n2715) );
  INV U3024 ( .A(n3202), .Y(n2716) );
  INV U3025 ( .A(n2716), .Y(n2717) );
  INV U3026 ( .A(n2521), .Y(n2718) );
  INV U3027 ( .A(n3837), .Y(n2719) );
  INV U3028 ( .A(n2719), .Y(n2720) );
  INV U3029 ( .A(n2520), .Y(n2721) );
  INV U3030 ( .A(n4992), .Y(n2722) );
  INV U3031 ( .A(n2722), .Y(disp1_sel[3]) );
  INV U3032 ( .A(\uut/mult_mant/shift_amount [5]), .Y(n2724) );
  INV U3033 ( .A(n2724), .Y(n2725) );
  INV U3034 ( .A(n4803), .Y(n2726) );
  INV U3035 ( .A(n2726), .Y(n2727) );
  INV U3036 ( .A(n4998), .Y(n2728) );
  INV U3037 ( .A(n2728), .Y(disp2_sel[3]) );
  INV U3038 ( .A(n4718), .Y(n2730) );
  INV U3039 ( .A(n2730), .Y(n2731) );
  INV U3040 ( .A(n4797), .Y(n2732) );
  INV U3041 ( .A(n2732), .Y(n2733) );
  INV U3042 ( .A(n3757), .Y(n2734) );
  INV U3043 ( .A(n2734), .Y(n2735) );
  INV U3044 ( .A(n5007), .Y(n2736) );
  INV U3045 ( .A(n2736), .Y(error) );
  INV U3046 ( .A(n2529), .Y(n2738) );
  INV U3047 ( .A(n2529), .Y(n2739) );
  INV U3048 ( .A(n4712), .Y(n2740) );
  INV U3049 ( .A(n2740), .Y(n2741) );
  INV U3050 ( .A(n4798), .Y(n2742) );
  INV U3051 ( .A(n2742), .Y(n2743) );
  INV U3052 ( .A(n2519), .Y(n2744) );
  INV U3053 ( .A(n2531), .Y(n2745) );
  INV U3054 ( .A(n2531), .Y(n2746) );
  INV U3055 ( .A(n3896), .Y(n2747) );
  INV U3056 ( .A(n2747), .Y(n2748) );
  INV U3057 ( .A(n3201), .Y(n2749) );
  INV U3058 ( .A(n2749), .Y(n2750) );
  INV U3059 ( .A(n3204), .Y(n2751) );
  INV U3060 ( .A(n2751), .Y(n2752) );
  INV U3061 ( .A(n4713), .Y(n2753) );
  INV U3062 ( .A(n2753), .Y(n2754) );
  INV U3063 ( .A(n2518), .Y(n2755) );
  INV U3064 ( .A(n3112), .Y(n2756) );
  INV U3065 ( .A(n3112), .Y(n2757) );
  INV U3066 ( .A(n2528), .Y(n2758) );
  INV U3067 ( .A(n2528), .Y(n2759) );
  INV U3068 ( .A(n2926), .Y(n2760) );
  INV U3069 ( .A(n2760), .Y(n2761) );
  INV U3070 ( .A(n3607), .Y(n2762) );
  INV U3071 ( .A(n2762), .Y(n2763) );
  INV U3072 ( .A(n2848), .Y(n2764) );
  INV U3073 ( .A(n2764), .Y(n2765) );
  INV U3074 ( .A(\uut/start ), .Y(n2766) );
  INV U3075 ( .A(\uut/start ), .Y(n2767) );
  INV U3076 ( .A(\uut/start ), .Y(n2768) );
  INV U3077 ( .A(n3446), .Y(n2769) );
  INV U3078 ( .A(n2769), .Y(n2770) );
  INV U3079 ( .A(n3436), .Y(n2771) );
  INV U3080 ( .A(n2771), .Y(n2772) );
  INV U3081 ( .A(n2739), .Y(n2773) );
  INV U3082 ( .A(n2738), .Y(n2774) );
  INV U3083 ( .A(n2739), .Y(n2775) );
  INV U3084 ( .A(n2738), .Y(n2776) );
  INV U3085 ( .A(n4161), .Y(n2777) );
  INV U3086 ( .A(n4161), .Y(n2778) );
  INV U3087 ( .A(n4161), .Y(n2779) );
  INV U3088 ( .A(n4161), .Y(n2780) );
  INV U3089 ( .A(n2779), .Y(n2781) );
  INV U3090 ( .A(n3471), .Y(n2782) );
  INV U3091 ( .A(n2782), .Y(n2783) );
  INV U3092 ( .A(input2_cnt[3]), .Y(n4786) );
  INV U3093 ( .A(input1_cnt[3]), .Y(n4871) );
  OAI2BB1 U3094 ( .A0N(n2528), .A1N(n2784), .B0(n2696), .Y(
        \uut/mult_mant/N299 ) );
  OAI2BB1 U3095 ( .A0N(n2697), .A1N(n2784), .B0(n2786), .Y(
        \uut/mult_mant/N298 ) );
  AOI21 U3096 ( .A0(n2787), .A1(\uut/start ), .B0(n2528), .Y(n2786) );
  NOR4BB U3097 ( .AN(ready), .BN(\uut/valid_q ), .C(error), .D(n2788), .Y(
        \uut/N66 ) );
  NAND3B U3098 ( .AN(\uut/mult_ready ), .B(n2789), .C(n2736), .Y(\uut/N64 ) );
  MX2 U3099 ( .A(\uut/exp_out[5] ), .B(\uut/exp_out[8] ), .S0(data_type), .Y(
        overflow) );
  MX2 U3100 ( .A(n2790), .B(n2791), .S0(n2541), .Y(n4880) );
  INV U3101 ( .A(n2792), .Y(n4881) );
  AOI21 U3102 ( .A0(\uut/exp_out[8] ), .A1(n2539), .B0(n2793), .Y(n2792) );
  MX2 U3103 ( .A(n2794), .B(n2795), .S0(n2796), .Y(n2793) );
  XNOR2 U3104 ( .A(n2797), .B(n2798), .Y(n2796) );
  ADDF U3105 ( .A(n2799), .B(n2800), .CI(n2801), .CO(n2798) );
  INV U3106 ( .A(n2802), .Y(n2800) );
  INV U3107 ( .A(n2803), .Y(n2799) );
  NOR2 U3108 ( .A(n2804), .B(n2805), .Y(n2797) );
  NOR2B U3109 ( .AN(n2806), .B(n2807), .Y(n2795) );
  OAI21 U3110 ( .A0(n2806), .A1(n2808), .B0(n2809), .Y(n2794) );
  OAI2BB1 U3111 ( .A0N(n2539), .A1N(\uut/exp_out[7] ), .B0(n2810), .Y(n4882)
         );
  MX2 U3112 ( .A(n2807), .B(n2809), .S0(n2806), .Y(n2810) );
  XNOR2 U3113 ( .A(n2804), .B(n2805), .Y(n2806) );
  AOI21 U3114 ( .A0(data_type), .A1(n2811), .B0(n2812), .Y(n2804) );
  NOR2B U3115 ( .AN(n2813), .B(n2814), .Y(n2809) );
  NOR2 U3116 ( .A(n2815), .B(n2808), .Y(n2814) );
  NAND2B U3117 ( .AN(n2808), .B(n2815), .Y(n2807) );
  NOR3B U3118 ( .AN(n2816), .B(n2817), .C(n2818), .Y(n2815) );
  OAI2BB1 U3119 ( .A0N(n2539), .A1N(\uut/exp_out[6] ), .B0(n2819), .Y(n4883)
         );
  AOI2BB1 U3120 ( .A0N(n2817), .A1N(n2820), .B0(n2821), .Y(n2819) );
  NOR4BB U3121 ( .AN(n2817), .BN(n2816), .C(n2818), .D(n2808), .Y(n2821) );
  NOR2B U3122 ( .AN(n2822), .B(n2823), .Y(n2820) );
  NOR2B U3123 ( .AN(n2818), .B(n2808), .Y(n2823) );
  ADDF U3124 ( .A(data_type), .B(n2812), .CI(n2811), .S(n2817) );
  AOI2BB2 U3125 ( .B0(n4961), .B1(n2824), .A0N(n2825), .A1N(n2826), .Y(n2812)
         );
  NOR2 U3126 ( .A(n4961), .B(n2824), .Y(n2826) );
  OAI2BB1 U3127 ( .A0N(n2539), .A1N(\uut/exp_out[5] ), .B0(n2827), .Y(n4884)
         );
  MX2 U3128 ( .A(n2822), .B(n2828), .S0(n2818), .Y(n2827) );
  ADDF U3129 ( .A(n2825), .B(n4961), .CI(n2824), .S(n2818) );
  AOI2BB1 U3130 ( .A0N(n2829), .A1N(n2830), .B0(n2831), .Y(n2825) );
  NAND2B U3131 ( .AN(n2808), .B(n2816), .Y(n2828) );
  NOR2B U3132 ( .AN(n2813), .B(n2832), .Y(n2822) );
  NOR2 U3133 ( .A(n2816), .B(n2808), .Y(n2832) );
  NOR3B U3134 ( .AN(n2833), .B(n2834), .C(n2835), .Y(n2816) );
  OAI2BB1 U3135 ( .A0N(n2539), .A1N(\uut/exp_out[4] ), .B0(n2836), .Y(n4885)
         );
  MX2 U3136 ( .A(n2837), .B(n2838), .S0(n2834), .Y(n2836) );
  MX2 U3137 ( .A(n2839), .B(n2840), .S0(n2830), .Y(n2834) );
  XNOR2 U3138 ( .A(data_type), .B(n2841), .Y(n2840) );
  NOR2 U3139 ( .A(n2829), .B(n2831), .Y(n2839) );
  NOR2 U3140 ( .A(n4961), .B(n2842), .Y(n2829) );
  OR2 U3141 ( .A(n2835), .B(n2843), .Y(n2838) );
  NOR2B U3142 ( .AN(n2844), .B(n2845), .Y(n2837) );
  NOR2B U3143 ( .AN(n2835), .B(n2808), .Y(n2845) );
  OAI2BB1 U3144 ( .A0N(\uut/in1_32_reg[0] ), .A1N(n2846), .B0(n2847), .Y(n4886) );
  AOI22 U3145 ( .A0(n2765), .A1(\uut/in1_16_reg[0] ), .B0(
        \uut/mult_mant/c1 [0]), .B1(n2767), .Y(n2847) );
  OAI2BB1 U3146 ( .A0N(\uut/in1_32_reg[1] ), .A1N(n2846), .B0(n2849), .Y(n4887) );
  AOI22 U3147 ( .A0(n2765), .A1(\uut/in1_16_reg[1] ), .B0(
        \uut/mult_mant/c1 [1]), .B1(n2766), .Y(n2849) );
  OAI2BB1 U3148 ( .A0N(\uut/in1_32_reg[2] ), .A1N(n2846), .B0(n2850), .Y(n4888) );
  AOI22 U3149 ( .A0(n2765), .A1(\uut/in1_16_reg[2] ), .B0(
        \uut/mult_mant/c1 [2]), .B1(n2768), .Y(n2850) );
  OAI2BB1 U3150 ( .A0N(\uut/in1_32_reg[3] ), .A1N(n2846), .B0(n2851), .Y(n4889) );
  AOI22 U3151 ( .A0(n2765), .A1(\uut/in1_16_reg[3] ), .B0(
        \uut/mult_mant/c1 [3]), .B1(n2767), .Y(n2851) );
  OAI2BB1 U3152 ( .A0N(\uut/in1_32_reg[4] ), .A1N(n2846), .B0(n2852), .Y(n4890) );
  AOI22 U3153 ( .A0(n2765), .A1(\uut/in1_16_reg[4] ), .B0(
        \uut/mult_mant/c1 [4]), .B1(n2766), .Y(n2852) );
  OAI2BB1 U3154 ( .A0N(\uut/in1_32_reg[5] ), .A1N(n2846), .B0(n2853), .Y(n4891) );
  AOI22 U3155 ( .A0(n2765), .A1(\uut/in1_16_reg[5] ), .B0(
        \uut/mult_mant/c1 [5]), .B1(n2768), .Y(n2853) );
  OAI2BB1 U3156 ( .A0N(\uut/in1_32_reg[6] ), .A1N(n2846), .B0(n2854), .Y(n4892) );
  AOI22 U3157 ( .A0(n2765), .A1(\uut/in1_16_reg[6] ), .B0(
        \uut/mult_mant/c1 [6]), .B1(n2767), .Y(n2854) );
  OAI2BB1 U3158 ( .A0N(\uut/in1_32_reg[7] ), .A1N(n2846), .B0(n2855), .Y(n4893) );
  AOI22 U3159 ( .A0(n2765), .A1(\uut/in1_16_reg[7] ), .B0(
        \uut/mult_mant/c1 [7]), .B1(n2766), .Y(n2855) );
  OAI2BB1 U3160 ( .A0N(\uut/in1_32_reg[8] ), .A1N(n2846), .B0(n2856), .Y(n4894) );
  AOI22 U3161 ( .A0(n2765), .A1(\uut/in1_16_reg[8] ), .B0(
        \uut/mult_mant/b1 [0]), .B1(n2768), .Y(n2856) );
  OAI2BB1 U3162 ( .A0N(\uut/in1_32_reg[9] ), .A1N(n2846), .B0(n2857), .Y(n4895) );
  AOI22 U3163 ( .A0(n2765), .A1(\uut/in1_16_reg[9] ), .B0(
        \uut/mult_mant/b1 [1]), .B1(n2767), .Y(n2857) );
  OAI21 U3164 ( .A0(n2533), .A1(n2764), .B0(n2859), .Y(n4896) );
  AOI22 U3165 ( .A0(n2846), .A1(\uut/in1_32_reg[10] ), .B0(
        \uut/mult_mant/b1 [2]), .B1(n2766), .Y(n2859) );
  OAI2BB1 U3166 ( .A0N(\uut/in2_32_reg[0] ), .A1N(n2846), .B0(n2860), .Y(n4897) );
  AOI22 U3167 ( .A0(n2765), .A1(\uut/in2_16_reg[0] ), .B0(
        \uut/mult_mant/c2 [0]), .B1(n2766), .Y(n2860) );
  OAI2BB1 U3168 ( .A0N(\uut/in2_32_reg[1] ), .A1N(n2846), .B0(n2861), .Y(n4898) );
  AOI22 U3169 ( .A0(n2765), .A1(\uut/in2_16_reg[1] ), .B0(
        \uut/mult_mant/c2 [1]), .B1(n2768), .Y(n2861) );
  OAI2BB1 U3170 ( .A0N(\uut/in2_32_reg[2] ), .A1N(n2846), .B0(n2862), .Y(n4899) );
  AOI22 U3171 ( .A0(n2765), .A1(\uut/in2_16_reg[2] ), .B0(
        \uut/mult_mant/c2 [2]), .B1(n2767), .Y(n2862) );
  OAI2BB1 U3172 ( .A0N(\uut/in2_32_reg[3] ), .A1N(n2846), .B0(n2863), .Y(n4900) );
  AOI22 U3173 ( .A0(n2765), .A1(\uut/in2_16_reg[3] ), .B0(
        \uut/mult_mant/c2 [3]), .B1(n2766), .Y(n2863) );
  OAI2BB1 U3174 ( .A0N(\uut/in2_32_reg[4] ), .A1N(n2846), .B0(n2864), .Y(n4901) );
  AOI22 U3175 ( .A0(n2765), .A1(\uut/in2_16_reg[4] ), .B0(
        \uut/mult_mant/c2 [4]), .B1(n2768), .Y(n2864) );
  OAI2BB1 U3176 ( .A0N(\uut/in2_32_reg[5] ), .A1N(n2846), .B0(n2865), .Y(n4902) );
  AOI22 U3177 ( .A0(n2765), .A1(\uut/in2_16_reg[5] ), .B0(
        \uut/mult_mant/c2 [5]), .B1(n2767), .Y(n2865) );
  OAI2BB1 U3178 ( .A0N(\uut/in2_32_reg[6] ), .A1N(n2846), .B0(n2866), .Y(n4903) );
  AOI22 U3179 ( .A0(n2765), .A1(\uut/in2_16_reg[6] ), .B0(
        \uut/mult_mant/c2 [6]), .B1(n2766), .Y(n2866) );
  OAI2BB1 U3180 ( .A0N(\uut/in2_32_reg[7] ), .A1N(n2846), .B0(n2867), .Y(n4904) );
  AOI22 U3181 ( .A0(n2765), .A1(\uut/in2_16_reg[7] ), .B0(
        \uut/mult_mant/c2 [7]), .B1(n2768), .Y(n2867) );
  OAI2BB1 U3182 ( .A0N(\uut/in2_32_reg[8] ), .A1N(n2846), .B0(n2868), .Y(n4905) );
  AOI22 U3183 ( .A0(n2765), .A1(\uut/in2_16_reg[8] ), .B0(
        \uut/mult_mant/b2 [0]), .B1(n2767), .Y(n2868) );
  OAI2BB1 U3184 ( .A0N(\uut/in2_32_reg[9] ), .A1N(n2846), .B0(n2869), .Y(n4906) );
  AOI22 U3185 ( .A0(n2765), .A1(\uut/in2_16_reg[9] ), .B0(
        \uut/mult_mant/b2 [1]), .B1(n2766), .Y(n2869) );
  OAI21 U3186 ( .A0(n2764), .A1(n2870), .B0(n2871), .Y(n4907) );
  AOI22 U3187 ( .A0(n2846), .A1(\uut/in2_32_reg[10] ), .B0(
        \uut/mult_mant/b2 [2]), .B1(n2768), .Y(n2871) );
  INV U3188 ( .A(n2544), .Y(n2846) );
  NOR2B U3189 ( .AN(\uut/start ), .B(data_type), .Y(n2848) );
  OAI21 U3190 ( .A0(n2872), .A1(n2808), .B0(n2873), .Y(n4908) );
  MX2 U3191 ( .A(n2874), .B(n2875), .S0(n2539), .Y(n2873) );
  INV U3192 ( .A(\uut/exp_out[0] ), .Y(n2875) );
  OAI2BB1 U3193 ( .A0N(n2876), .A1N(n2877), .B0(n2878), .Y(n2874) );
  OAI2BB1 U3194 ( .A0N(n2539), .A1N(\uut/exp_out[3] ), .B0(n2879), .Y(n4909)
         );
  MX2 U3195 ( .A(n2844), .B(n2843), .S0(n2835), .Y(n2879) );
  XNOR2 U3196 ( .A(n2880), .B(n2881), .Y(n2835) );
  NAND2B U3197 ( .AN(n2808), .B(n2833), .Y(n2843) );
  NOR2B U3198 ( .AN(n2813), .B(n2882), .Y(n2844) );
  NOR2 U3199 ( .A(n2833), .B(n2808), .Y(n2882) );
  NOR2B U3200 ( .AN(n2883), .B(n2884), .Y(n2833) );
  INV U3201 ( .A(n2885), .Y(n4910) );
  AOI21 U3202 ( .A0(n2539), .A1(\uut/exp_out[2] ), .B0(n2886), .Y(n2885) );
  MX2 U3203 ( .A(n2887), .B(n2888), .S0(n2884), .Y(n2886) );
  XOR2 U3204 ( .A(n2889), .B(n2890), .Y(n2884) );
  NOR2B U3205 ( .AN(n2883), .B(n2808), .Y(n2888) );
  OAI21 U3206 ( .A0(n2883), .A1(n2808), .B0(n2813), .Y(n2887) );
  OAI222 U3207 ( .A0(n2891), .A1(n2538), .B0(n2813), .B1(n2892), .C0(n2808), 
        .C1(n2893), .Y(n4911) );
  NAND2B U3208 ( .AN(n2539), .B(\uut/normalize ), .Y(n2808) );
  AOI2BB1 U3209 ( .A0N(n2893), .A1N(n2872), .B0(n2883), .Y(n2892) );
  NOR2B U3210 ( .AN(n2893), .B(n2876), .Y(n2883) );
  INV U3211 ( .A(n2872), .Y(n2876) );
  OR2 U3212 ( .A(n2539), .B(\uut/normalize ), .Y(n2813) );
  INV U3213 ( .A(\uut/exp_out[1] ), .Y(n2891) );
  OAI211 U3214 ( .A0(enter), .A1(n2538), .B0(n2877), .C0(n2878), .Y(n4912) );
  NAND2B U3215 ( .AN(n2805), .B(n2894), .Y(n2877) );
  NOR4BB U3216 ( .AN(n2895), .BN(\uut/more_than_1 ), .C(n2896), .D(n2897), .Y(
        n2894) );
  MX2 U3217 ( .A(data_type), .B(n2811), .S0(n2824), .Y(n2897) );
  ADDF U3218 ( .A(n2898), .B(n2899), .CI(n2900), .S(n2824) );
  INV U3219 ( .A(n2901), .Y(n2811) );
  XOR2 U3220 ( .A(n2533), .B(n2902), .Y(n2896) );
  AOI211 U3221 ( .A0(n2841), .A1(n2901), .B0(n2831), .C0(n2830), .Y(n2895) );
  NAND2 U3222 ( .A(n2880), .B(n2881), .Y(n2830) );
  ADDF U3223 ( .A(n2903), .B(n2904), .CI(n2905), .S(n2881) );
  INV U3224 ( .A(n2906), .Y(n2904) );
  INV U3225 ( .A(n2907), .Y(n2903) );
  NOR2B U3226 ( .AN(n2890), .B(n2889), .Y(n2880) );
  ADDF U3227 ( .A(n2908), .B(n2909), .CI(n2910), .S(n2889) );
  INV U3228 ( .A(n2911), .Y(n2908) );
  NOR2B U3229 ( .AN(n2893), .B(n2872), .Y(n2890) );
  XNOR2 U3230 ( .A(n2912), .B(n2913), .Y(n2872) );
  ADDF U3231 ( .A(n2914), .B(n2915), .CI(n2916), .S(n2893) );
  NOR2B U3232 ( .AN(n2842), .B(data_type), .Y(n2831) );
  INV U3233 ( .A(n2841), .Y(n2842) );
  ADDF U3234 ( .A(n2917), .B(n2918), .CI(n2919), .S(n2901) );
  ADDF U3235 ( .A(n2920), .B(n2921), .CI(n2922), .S(n2841) );
  INV U3236 ( .A(n2923), .Y(n2920) );
  ADDF U3237 ( .A(n2803), .B(n2802), .CI(n2801), .S(n2805) );
  ADDF U3238 ( .A(n2917), .B(n2918), .CI(n2919), .CO(n2801) );
  ADDF U3239 ( .A(n2898), .B(n2899), .CI(n2900), .CO(n2919) );
  ADDF U3240 ( .A(n2923), .B(n2921), .CI(n2922), .CO(n2900) );
  MX2 U3241 ( .A(\uut/in2_16_reg[14] ), .B(\uut/in2_32_reg[27] ), .S0(
        data_type), .Y(n2921) );
  ADDF U3242 ( .A(n2905), .B(n2907), .CI(n2906), .CO(n2923) );
  MX2 U3243 ( .A(\uut/in2_16_reg[13] ), .B(\uut/in2_32_reg[26] ), .S0(
        data_type), .Y(n2906) );
  ADDF U3244 ( .A(n2909), .B(n2911), .CI(n2910), .CO(n2905) );
  MX2 U3245 ( .A(\uut/in2_16_reg[12] ), .B(\uut/in2_32_reg[25] ), .S0(
        data_type), .Y(n2910) );
  ADDF U3246 ( .A(n2914), .B(n2915), .CI(n2916), .CO(n2909) );
  MX2 U3247 ( .A(\uut/in2_16_reg[11] ), .B(\uut/in2_32_reg[24] ), .S0(
        data_type), .Y(n2916) );
  NOR2B U3248 ( .AN(n2913), .B(n2924), .Y(n2914) );
  MX2 U3249 ( .A(\uut/in2_16_reg[10] ), .B(\uut/in2_32_reg[23] ), .S0(
        data_type), .Y(n2913) );
  NOR2B U3250 ( .AN(\uut/in2_32_reg[28] ), .B(n4961), .Y(n2899) );
  NOR2B U3251 ( .AN(\uut/in2_32_reg[29] ), .B(n4961), .Y(n2918) );
  OAI222 U3252 ( .A0(n2925), .A1(n2926), .B0(n2759), .B1(n2927), .C0(n2757), 
        .C1(n2928), .Y(n4913) );
  ADDF U3253 ( .A(n2929), .B(\uut/mult_mant/temp_product[45] ), .CI(n2930), 
        .S(n2927) );
  OAI222 U3254 ( .A0(n2761), .A1(n2928), .B0(n2758), .B1(n2931), .C0(n2932), 
        .C1(n2756), .Y(n4914) );
  ADDF U3255 ( .A(\uut/mult_mant/temp_product[44] ), .B(n2933), .CI(n2934), 
        .S(n2931) );
  OAI222 U3256 ( .A0(n2761), .A1(n2932), .B0(n2759), .B1(n2935), .C0(n2936), 
        .C1(n2757), .Y(n4915) );
  ADDF U3257 ( .A(\uut/mult_mant/temp_product[43] ), .B(n2937), .CI(n2938), 
        .S(n2935) );
  OAI222 U3258 ( .A0(n2761), .A1(n2936), .B0(n2758), .B1(n2939), .C0(n2940), 
        .C1(n2756), .Y(n4916) );
  ADDF U3259 ( .A(\uut/mult_mant/temp_product[42] ), .B(n2941), .CI(n2942), 
        .S(n2939) );
  OAI222 U3260 ( .A0(n2926), .A1(n2940), .B0(n2759), .B1(n2943), .C0(n2944), 
        .C1(n2757), .Y(n4917) );
  ADDF U3261 ( .A(\uut/mult_mant/temp_product[41] ), .B(n2945), .CI(n2946), 
        .S(n2943) );
  OAI222 U3262 ( .A0(n2761), .A1(n2944), .B0(n2758), .B1(n2947), .C0(n2948), 
        .C1(n2756), .Y(n4918) );
  ADDF U3263 ( .A(\uut/mult_mant/temp_product[40] ), .B(n2949), .CI(n2950), 
        .S(n2947) );
  OAI222 U3264 ( .A0(n2926), .A1(n2948), .B0(n2951), .B1(n2759), .C0(n2757), 
        .C1(n2952), .Y(n4919) );
  ADDF U3265 ( .A(n2953), .B(\uut/mult_mant/temp_product[39] ), .CI(n2954), 
        .S(n2951) );
  OAI222 U3266 ( .A0(n2761), .A1(n2952), .B0(n2955), .B1(n2758), .C0(n2756), 
        .C1(n2956), .Y(n4920) );
  ADDF U3267 ( .A(n2957), .B(\uut/mult_mant/temp_product[38] ), .CI(n2958), 
        .S(n2955) );
  OAI222 U3268 ( .A0(n2926), .A1(n2956), .B0(n2959), .B1(n2759), .C0(n2757), 
        .C1(n2960), .Y(n4921) );
  ADDF U3269 ( .A(n2961), .B(\uut/mult_mant/temp_product[37] ), .CI(n2962), 
        .S(n2959) );
  OAI222 U3270 ( .A0(n2761), .A1(n2960), .B0(n2963), .B1(n2758), .C0(n2756), 
        .C1(n2964), .Y(n4922) );
  ADDF U3271 ( .A(n2965), .B(\uut/mult_mant/temp_product[36] ), .CI(n2966), 
        .S(n2963) );
  OAI222 U3272 ( .A0(n2926), .A1(n2964), .B0(n2967), .B1(n2759), .C0(n2757), 
        .C1(n2968), .Y(n4923) );
  ADDF U3273 ( .A(n2969), .B(\uut/mult_mant/temp_product[35] ), .CI(n2970), 
        .S(n2967) );
  OAI222 U3274 ( .A0(n2761), .A1(n2968), .B0(n2971), .B1(n2758), .C0(n2756), 
        .C1(n2972), .Y(n4924) );
  ADDF U3275 ( .A(n2973), .B(\uut/mult_mant/temp_product[34] ), .CI(n2974), 
        .S(n2971) );
  OAI222 U3276 ( .A0(n2926), .A1(n2972), .B0(n2975), .B1(n2759), .C0(n2757), 
        .C1(n2976), .Y(n4925) );
  ADDF U3277 ( .A(n2977), .B(\uut/mult_mant/temp_product[33] ), .CI(n2978), 
        .S(n2975) );
  OAI222 U3278 ( .A0(n2761), .A1(n2976), .B0(n2979), .B1(n2758), .C0(n2756), 
        .C1(n2980), .Y(n4926) );
  ADDF U3279 ( .A(n2981), .B(\uut/mult_mant/temp_product[32] ), .CI(n2982), 
        .S(n2979) );
  OAI222 U3280 ( .A0(n2926), .A1(n2980), .B0(n2983), .B1(n2759), .C0(n2757), 
        .C1(n2984), .Y(n4927) );
  ADDF U3281 ( .A(n2985), .B(\uut/mult_mant/temp_product[31] ), .CI(n2986), 
        .S(n2983) );
  OAI222 U3282 ( .A0(n2761), .A1(n2984), .B0(n2987), .B1(n2758), .C0(n2756), 
        .C1(n2988), .Y(n4928) );
  ADDF U3283 ( .A(n2989), .B(\uut/mult_mant/temp_product[30] ), .CI(n2990), 
        .S(n2987) );
  OAI222 U3284 ( .A0(n2926), .A1(n2988), .B0(n2991), .B1(n2759), .C0(n2757), 
        .C1(n2992), .Y(n4929) );
  ADDF U3285 ( .A(n2993), .B(\uut/mult_mant/temp_product[29] ), .CI(n2994), 
        .S(n2991) );
  OAI222 U3286 ( .A0(n2761), .A1(n2992), .B0(n2995), .B1(n2758), .C0(n2756), 
        .C1(n2996), .Y(n4930) );
  ADDF U3287 ( .A(n2997), .B(\uut/mult_mant/temp_product[28] ), .CI(n2998), 
        .S(n2995) );
  OAI222 U3288 ( .A0(n2926), .A1(n2996), .B0(n2999), .B1(n2759), .C0(n2757), 
        .C1(n3000), .Y(n4931) );
  ADDF U3289 ( .A(n3001), .B(\uut/mult_mant/temp_product[27] ), .CI(n3002), 
        .S(n2999) );
  OAI222 U3290 ( .A0(n2761), .A1(n3000), .B0(n3003), .B1(n2758), .C0(n2756), 
        .C1(n3004), .Y(n4932) );
  ADDF U3291 ( .A(n3005), .B(\uut/mult_mant/temp_product[26] ), .CI(n3006), 
        .S(n3003) );
  OAI222 U3292 ( .A0(n2926), .A1(n3004), .B0(n3007), .B1(n2759), .C0(n2757), 
        .C1(n3008), .Y(n4933) );
  ADDF U3293 ( .A(n3009), .B(\uut/mult_mant/temp_product[25] ), .CI(n3010), 
        .S(n3007) );
  OAI222 U3294 ( .A0(n2761), .A1(n3008), .B0(n3011), .B1(n2758), .C0(n2756), 
        .C1(n3012), .Y(n4934) );
  ADDF U3295 ( .A(n3013), .B(\uut/mult_mant/temp_product[24] ), .CI(n3014), 
        .S(n3011) );
  OAI222 U3296 ( .A0(n2926), .A1(n3012), .B0(n3015), .B1(n2759), .C0(n2757), 
        .C1(n3016), .Y(n4935) );
  ADDF U3297 ( .A(n3017), .B(\uut/mult_mant/temp_product[23] ), .CI(n3018), 
        .S(n3015) );
  OAI222 U3298 ( .A0(n2761), .A1(n3016), .B0(n3019), .B1(n2758), .C0(n2756), 
        .C1(n3020), .Y(n4936) );
  ADDF U3299 ( .A(n3021), .B(\uut/mult_mant/temp_product[22] ), .CI(n3022), 
        .S(n3019) );
  OAI222 U3300 ( .A0(n2926), .A1(n3020), .B0(n3023), .B1(n2759), .C0(n2757), 
        .C1(n3024), .Y(n4937) );
  ADDF U3301 ( .A(n3025), .B(\uut/mult_mant/temp_product[21] ), .CI(n3026), 
        .S(n3023) );
  INV U3302 ( .A(\uut/mult_mant/temp_product[22] ), .Y(n3020) );
  OAI222 U3303 ( .A0(n2761), .A1(n3024), .B0(n3027), .B1(n2758), .C0(n2756), 
        .C1(n3028), .Y(n4938) );
  ADDF U3304 ( .A(n3029), .B(\uut/mult_mant/temp_product[20] ), .CI(n3030), 
        .S(n3027) );
  INV U3305 ( .A(\uut/mult_mant/temp_product[21] ), .Y(n3024) );
  OAI222 U3306 ( .A0(n2926), .A1(n3028), .B0(n3031), .B1(n2759), .C0(n2757), 
        .C1(n3032), .Y(n4939) );
  ADDF U3307 ( .A(n3033), .B(\uut/mult_mant/temp_product[19] ), .CI(n3034), 
        .S(n3031) );
  INV U3308 ( .A(\uut/mult_mant/temp_product[20] ), .Y(n3028) );
  OAI222 U3309 ( .A0(n2761), .A1(n3032), .B0(n3035), .B1(n2758), .C0(n2756), 
        .C1(n3036), .Y(n4940) );
  ADDF U3310 ( .A(n3037), .B(\uut/mult_mant/temp_product[18] ), .CI(n3038), 
        .S(n3035) );
  OAI222 U3311 ( .A0(n2926), .A1(n3036), .B0(n3039), .B1(n2759), .C0(n2757), 
        .C1(n3040), .Y(n4941) );
  ADDF U3312 ( .A(n3041), .B(\uut/mult_mant/temp_product[17] ), .CI(n3042), 
        .S(n3039) );
  OAI222 U3313 ( .A0(n2761), .A1(n3040), .B0(n3043), .B1(n2758), .C0(n2756), 
        .C1(n3044), .Y(n4942) );
  ADDF U3314 ( .A(n3045), .B(\uut/mult_mant/temp_product[16] ), .CI(n3046), 
        .S(n3043) );
  OAI222 U3315 ( .A0(n2926), .A1(n3044), .B0(n2759), .B1(n3047), .C0(n3048), 
        .C1(n2757), .Y(n4943) );
  ADDF U3316 ( .A(\uut/mult_mant/temp_product[15] ), .B(n3049), .CI(n3050), 
        .S(n3047) );
  OAI222 U3317 ( .A0(n2761), .A1(n3048), .B0(n2758), .B1(n3051), .C0(n3052), 
        .C1(n2756), .Y(n4944) );
  ADDF U3318 ( .A(\uut/mult_mant/temp_product[14] ), .B(n3053), .CI(n3054), 
        .S(n3051) );
  OAI222 U3319 ( .A0(n2926), .A1(n3052), .B0(n2759), .B1(n3055), .C0(n3056), 
        .C1(n2757), .Y(n4945) );
  ADDF U3320 ( .A(\uut/mult_mant/temp_product[13] ), .B(n3057), .CI(n3058), 
        .S(n3055) );
  OAI222 U3321 ( .A0(n2761), .A1(n3056), .B0(n2758), .B1(n3059), .C0(n3060), 
        .C1(n2756), .Y(n4946) );
  ADDF U3322 ( .A(\uut/mult_mant/temp_product[12] ), .B(n3061), .CI(n3062), 
        .S(n3059) );
  OAI222 U3323 ( .A0(n2926), .A1(n3060), .B0(n2759), .B1(n3063), .C0(n3064), 
        .C1(n2757), .Y(n4947) );
  ADDF U3324 ( .A(\uut/mult_mant/temp_product[11] ), .B(n3065), .CI(n3066), 
        .S(n3063) );
  OAI222 U3325 ( .A0(n2761), .A1(n3064), .B0(n2758), .B1(n3067), .C0(n3068), 
        .C1(n2756), .Y(n4948) );
  ADDF U3326 ( .A(\uut/mult_mant/temp_product[10] ), .B(n3069), .CI(n3070), 
        .S(n3067) );
  OAI222 U3327 ( .A0(n2926), .A1(n3068), .B0(n2759), .B1(n3071), .C0(n3072), 
        .C1(n2757), .Y(n4949) );
  ADDF U3328 ( .A(\uut/mult_mant/temp_product[9] ), .B(n3073), .CI(n3074), .S(
        n3071) );
  OAI222 U3329 ( .A0(n2761), .A1(n3072), .B0(n2758), .B1(n3075), .C0(n3076), 
        .C1(n2756), .Y(n4950) );
  ADDF U3330 ( .A(\uut/mult_mant/temp_product[8] ), .B(n3077), .CI(n3078), .S(
        n3075) );
  INV U3331 ( .A(\uut/mult_mant/temp_product[9] ), .Y(n3072) );
  OAI222 U3332 ( .A0(n2926), .A1(n3076), .B0(n2759), .B1(n3079), .C0(n3080), 
        .C1(n2757), .Y(n4951) );
  ADDF U3333 ( .A(\uut/mult_mant/temp_product[7] ), .B(n3081), .CI(n3082), .S(
        n3079) );
  INV U3334 ( .A(\uut/mult_mant/temp_product[8] ), .Y(n3076) );
  OAI222 U3335 ( .A0(n2761), .A1(n3080), .B0(n2758), .B1(n3083), .C0(n3084), 
        .C1(n2756), .Y(n4952) );
  ADDF U3336 ( .A(\uut/mult_mant/temp_product[6] ), .B(n3085), .CI(n3086), .S(
        n3083) );
  INV U3337 ( .A(\uut/mult_mant/temp_product[7] ), .Y(n3080) );
  OAI222 U3338 ( .A0(n2926), .A1(n3084), .B0(n2759), .B1(n3087), .C0(n3088), 
        .C1(n2757), .Y(n4953) );
  ADDF U3339 ( .A(\uut/mult_mant/temp_product[5] ), .B(n3089), .CI(n3090), .S(
        n3087) );
  INV U3340 ( .A(\uut/mult_mant/temp_product[6] ), .Y(n3084) );
  OAI222 U3341 ( .A0(n2761), .A1(n3088), .B0(n2758), .B1(n3091), .C0(n3092), 
        .C1(n2756), .Y(n4954) );
  ADDF U3342 ( .A(\uut/mult_mant/temp_product[4] ), .B(n3093), .CI(n3094), .S(
        n3091) );
  INV U3343 ( .A(\uut/mult_mant/temp_product[5] ), .Y(n3088) );
  OAI222 U3344 ( .A0(n2926), .A1(n3092), .B0(n2759), .B1(n3095), .C0(n3096), 
        .C1(n2757), .Y(n4955) );
  ADDF U3345 ( .A(n3097), .B(n3098), .CI(\uut/mult_mant/temp_product[3] ), .S(
        n3095) );
  INV U3346 ( .A(\uut/mult_mant/temp_product[4] ), .Y(n3092) );
  OAI222 U3347 ( .A0(n2761), .A1(n3096), .B0(n2758), .B1(n3099), .C0(n3100), 
        .C1(n2756), .Y(n4956) );
  ADDF U3348 ( .A(\uut/mult_mant/temp_product[2] ), .B(n3101), .CI(n3102), .S(
        n3099) );
  INV U3349 ( .A(\uut/mult_mant/temp_product[3] ), .Y(n3096) );
  OAI222 U3350 ( .A0(n2926), .A1(n3100), .B0(n3103), .B1(n2759), .C0(n2757), 
        .C1(n3104), .Y(n4957) );
  ADDF U3351 ( .A(n3105), .B(\uut/mult_mant/temp_product[1] ), .CI(n3106), .S(
        n3103) );
  INV U3352 ( .A(\uut/mult_mant/temp_product[2] ), .Y(n3100) );
  OAI222 U3353 ( .A0(n2761), .A1(n3104), .B0(n3107), .B1(n2758), .C0(n2756), 
        .C1(n3108), .Y(n4958) );
  INV U3354 ( .A(\uut/mult_mant/temp_product[0] ), .Y(n3108) );
  XNOR2 U3355 ( .A(n3109), .B(\uut/mult_mant/temp_product[0] ), .Y(n3107) );
  INV U3356 ( .A(\uut/mult_mant/temp_product[1] ), .Y(n3104) );
  OAI222 U3357 ( .A0(n2925), .A1(n2757), .B0(n2759), .B1(n3110), .C0(n3111), 
        .C1(n2926), .Y(n4959) );
  NAND2B U3358 ( .AN(n3112), .B(n2641), .Y(n2926) );
  ADDF U3359 ( .A(\uut/mult_mant/temp_product[46] ), .B(n3113), .CI(n3114), 
        .S(n3110) );
  OAI2BB2 U3360 ( .B0(n3111), .B1(n2756), .A0N(n2528), .A1N(n3115), .Y(n4960)
         );
  ADDF U3361 ( .A(\uut/mult_mant/temp_product[47] ), .B(n3116), .CI(n3117), 
        .S(n3115) );
  OAI22 U3362 ( .A0(n3113), .A1(n2925), .B0(n3118), .B1(n3119), .Y(n3117) );
  INV U3363 ( .A(n3114), .Y(n3119) );
  NOR2B U3364 ( .AN(n3120), .B(n2724), .Y(n3114) );
  NOR2B U3365 ( .AN(n3113), .B(\uut/mult_mant/temp_product[46] ), .Y(n3118) );
  INV U3366 ( .A(\uut/mult_mant/temp_product[46] ), .Y(n2925) );
  AOI2BB2 U3367 ( .B0(\uut/mult_mant/temp_product[45] ), .B1(n3121), .A0N(
        n3122), .A1N(n3123), .Y(n3113) );
  INV U3368 ( .A(n2930), .Y(n3123) );
  NOR2B U3369 ( .AN(n3124), .B(n2724), .Y(n2930) );
  NOR2B U3370 ( .AN(n2929), .B(\uut/mult_mant/temp_product[45] ), .Y(n3122) );
  INV U3371 ( .A(n2929), .Y(n3121) );
  AOI2BB2 U3372 ( .B0(\uut/mult_mant/temp_product[44] ), .B1(n2933), .A0N(
        n3125), .A1N(n2934), .Y(n2929) );
  NAND2 U3373 ( .A(n2725), .B(n3126), .Y(n2934) );
  NOR2 U3374 ( .A(\uut/mult_mant/temp_product[44] ), .B(n2933), .Y(n3125) );
  OAI2BB2 U3375 ( .B0(n3127), .B1(n2938), .A0N(
        \uut/mult_mant/temp_product[43] ), .A1N(n2937), .Y(n2933) );
  NAND2 U3376 ( .A(n2725), .B(n3128), .Y(n2938) );
  NOR2 U3377 ( .A(\uut/mult_mant/temp_product[43] ), .B(n2937), .Y(n3127) );
  OAI2BB2 U3378 ( .B0(n3129), .B1(n2942), .A0N(
        \uut/mult_mant/temp_product[42] ), .A1N(n2941), .Y(n2937) );
  NAND2 U3379 ( .A(n2725), .B(n3130), .Y(n2942) );
  NOR2 U3380 ( .A(\uut/mult_mant/temp_product[42] ), .B(n2941), .Y(n3129) );
  OAI2BB2 U3381 ( .B0(n3131), .B1(n2946), .A0N(
        \uut/mult_mant/temp_product[41] ), .A1N(n2945), .Y(n2941) );
  NAND2 U3382 ( .A(n2725), .B(n3132), .Y(n2946) );
  NOR2 U3383 ( .A(\uut/mult_mant/temp_product[41] ), .B(n2945), .Y(n3131) );
  OAI2BB2 U3384 ( .B0(n3133), .B1(n2950), .A0N(
        \uut/mult_mant/temp_product[40] ), .A1N(n2949), .Y(n2945) );
  NAND2 U3385 ( .A(n2725), .B(n3134), .Y(n2950) );
  NOR2 U3386 ( .A(\uut/mult_mant/temp_product[40] ), .B(n2949), .Y(n3133) );
  OAI2BB2 U3387 ( .B0(n2953), .B1(n3135), .A0N(
        \uut/mult_mant/temp_product[39] ), .A1N(n2954), .Y(n2949) );
  NOR2 U3388 ( .A(\uut/mult_mant/temp_product[39] ), .B(n2954), .Y(n3135) );
  OAI2BB2 U3389 ( .B0(n2957), .B1(n3136), .A0N(
        \uut/mult_mant/temp_product[38] ), .A1N(n2958), .Y(n2954) );
  NOR2 U3390 ( .A(\uut/mult_mant/temp_product[38] ), .B(n2958), .Y(n3136) );
  OAI2BB2 U3391 ( .B0(n2961), .B1(n3137), .A0N(
        \uut/mult_mant/temp_product[37] ), .A1N(n2962), .Y(n2958) );
  NOR2 U3392 ( .A(\uut/mult_mant/temp_product[37] ), .B(n2962), .Y(n3137) );
  OAI2BB2 U3393 ( .B0(n2965), .B1(n3138), .A0N(
        \uut/mult_mant/temp_product[36] ), .A1N(n2966), .Y(n2962) );
  NOR2 U3394 ( .A(\uut/mult_mant/temp_product[36] ), .B(n2966), .Y(n3138) );
  OAI2BB2 U3395 ( .B0(n2969), .B1(n3139), .A0N(
        \uut/mult_mant/temp_product[35] ), .A1N(n2970), .Y(n2966) );
  NOR2 U3396 ( .A(\uut/mult_mant/temp_product[35] ), .B(n2970), .Y(n3139) );
  OAI2BB2 U3397 ( .B0(n2973), .B1(n3140), .A0N(
        \uut/mult_mant/temp_product[34] ), .A1N(n2974), .Y(n2970) );
  NOR2 U3398 ( .A(\uut/mult_mant/temp_product[34] ), .B(n2974), .Y(n3140) );
  OAI2BB2 U3399 ( .B0(n2977), .B1(n3141), .A0N(
        \uut/mult_mant/temp_product[33] ), .A1N(n2978), .Y(n2974) );
  NOR2 U3400 ( .A(\uut/mult_mant/temp_product[33] ), .B(n2978), .Y(n3141) );
  OAI2BB2 U3401 ( .B0(n2981), .B1(n3142), .A0N(
        \uut/mult_mant/temp_product[32] ), .A1N(n2982), .Y(n2978) );
  NOR2 U3402 ( .A(\uut/mult_mant/temp_product[32] ), .B(n2982), .Y(n3142) );
  OAI2BB2 U3403 ( .B0(n2985), .B1(n3143), .A0N(
        \uut/mult_mant/temp_product[31] ), .A1N(n2986), .Y(n2982) );
  NOR2 U3404 ( .A(\uut/mult_mant/temp_product[31] ), .B(n2986), .Y(n3143) );
  OAI2BB2 U3405 ( .B0(n2989), .B1(n3144), .A0N(
        \uut/mult_mant/temp_product[30] ), .A1N(n2990), .Y(n2986) );
  NOR2 U3406 ( .A(\uut/mult_mant/temp_product[30] ), .B(n2990), .Y(n3144) );
  OAI2BB2 U3407 ( .B0(n2993), .B1(n3145), .A0N(
        \uut/mult_mant/temp_product[29] ), .A1N(n2994), .Y(n2990) );
  NOR2 U3408 ( .A(\uut/mult_mant/temp_product[29] ), .B(n2994), .Y(n3145) );
  OAI2BB2 U3409 ( .B0(n2997), .B1(n3146), .A0N(
        \uut/mult_mant/temp_product[28] ), .A1N(n2998), .Y(n2994) );
  NOR2 U3410 ( .A(\uut/mult_mant/temp_product[28] ), .B(n2998), .Y(n3146) );
  OAI2BB2 U3411 ( .B0(n3001), .B1(n3147), .A0N(
        \uut/mult_mant/temp_product[27] ), .A1N(n3002), .Y(n2998) );
  NOR2 U3412 ( .A(\uut/mult_mant/temp_product[27] ), .B(n3002), .Y(n3147) );
  OAI2BB2 U3413 ( .B0(n3005), .B1(n3148), .A0N(
        \uut/mult_mant/temp_product[26] ), .A1N(n3006), .Y(n3002) );
  NOR2 U3414 ( .A(\uut/mult_mant/temp_product[26] ), .B(n3006), .Y(n3148) );
  OAI2BB2 U3415 ( .B0(n3009), .B1(n3149), .A0N(
        \uut/mult_mant/temp_product[25] ), .A1N(n3010), .Y(n3006) );
  NOR2 U3416 ( .A(\uut/mult_mant/temp_product[25] ), .B(n3010), .Y(n3149) );
  OAI2BB2 U3417 ( .B0(n3013), .B1(n3150), .A0N(
        \uut/mult_mant/temp_product[24] ), .A1N(n3014), .Y(n3010) );
  NOR2 U3418 ( .A(\uut/mult_mant/temp_product[24] ), .B(n3014), .Y(n3150) );
  OAI2BB2 U3419 ( .B0(n3017), .B1(n3151), .A0N(
        \uut/mult_mant/temp_product[23] ), .A1N(n3018), .Y(n3014) );
  NOR2 U3420 ( .A(\uut/mult_mant/temp_product[23] ), .B(n3018), .Y(n3151) );
  OAI2BB2 U3421 ( .B0(n3021), .B1(n3152), .A0N(
        \uut/mult_mant/temp_product[22] ), .A1N(n3022), .Y(n3018) );
  NOR2 U3422 ( .A(\uut/mult_mant/temp_product[22] ), .B(n3022), .Y(n3152) );
  OAI2BB2 U3423 ( .B0(n3025), .B1(n3153), .A0N(
        \uut/mult_mant/temp_product[21] ), .A1N(n3026), .Y(n3022) );
  NOR2 U3424 ( .A(\uut/mult_mant/temp_product[21] ), .B(n3026), .Y(n3153) );
  OAI2BB2 U3425 ( .B0(n3029), .B1(n3154), .A0N(
        \uut/mult_mant/temp_product[20] ), .A1N(n3030), .Y(n3026) );
  NOR2 U3426 ( .A(\uut/mult_mant/temp_product[20] ), .B(n3030), .Y(n3154) );
  OAI2BB2 U3427 ( .B0(n3033), .B1(n3155), .A0N(
        \uut/mult_mant/temp_product[19] ), .A1N(n3034), .Y(n3030) );
  NOR2 U3428 ( .A(\uut/mult_mant/temp_product[19] ), .B(n3034), .Y(n3155) );
  OAI2BB2 U3429 ( .B0(n3037), .B1(n3156), .A0N(
        \uut/mult_mant/temp_product[18] ), .A1N(n3038), .Y(n3034) );
  NOR2 U3430 ( .A(\uut/mult_mant/temp_product[18] ), .B(n3038), .Y(n3156) );
  OAI2BB2 U3431 ( .B0(n3041), .B1(n3157), .A0N(
        \uut/mult_mant/temp_product[17] ), .A1N(n3042), .Y(n3038) );
  NOR2 U3432 ( .A(\uut/mult_mant/temp_product[17] ), .B(n3042), .Y(n3157) );
  OAI2BB2 U3433 ( .B0(n3045), .B1(n3158), .A0N(
        \uut/mult_mant/temp_product[16] ), .A1N(n3046), .Y(n3042) );
  NOR2 U3434 ( .A(\uut/mult_mant/temp_product[16] ), .B(n3046), .Y(n3158) );
  OAI2BB2 U3435 ( .B0(n3159), .B1(n3050), .A0N(
        \uut/mult_mant/temp_product[15] ), .A1N(n3049), .Y(n3046) );
  OR2 U3436 ( .A(n2725), .B(n3160), .Y(n3050) );
  NOR2 U3437 ( .A(\uut/mult_mant/temp_product[15] ), .B(n3049), .Y(n3159) );
  OAI2BB2 U3438 ( .B0(n3161), .B1(n3054), .A0N(
        \uut/mult_mant/temp_product[14] ), .A1N(n3053), .Y(n3049) );
  NAND2B U3439 ( .AN(n2725), .B(n3120), .Y(n3054) );
  NOR2B U3440 ( .AN(n3162), .B(n2549), .Y(n3120) );
  MX2 U3441 ( .A(n3163), .B(n3164), .S0(n2699), .Y(n3162) );
  NOR2 U3442 ( .A(\uut/mult_mant/temp_product[14] ), .B(n3053), .Y(n3161) );
  OAI2BB2 U3443 ( .B0(n3165), .B1(n3058), .A0N(
        \uut/mult_mant/temp_product[13] ), .A1N(n3057), .Y(n3053) );
  NAND2B U3444 ( .AN(n2725), .B(n3124), .Y(n3058) );
  NOR2B U3445 ( .AN(n3166), .B(n2549), .Y(n3124) );
  MX2 U3446 ( .A(n3167), .B(n3168), .S0(n2699), .Y(n3166) );
  NOR2 U3447 ( .A(\uut/mult_mant/temp_product[13] ), .B(n3057), .Y(n3165) );
  OAI2BB2 U3448 ( .B0(n3169), .B1(n3062), .A0N(
        \uut/mult_mant/temp_product[12] ), .A1N(n3061), .Y(n3057) );
  NAND2B U3449 ( .AN(n2725), .B(n3126), .Y(n3062) );
  NOR2B U3450 ( .AN(n3170), .B(n2549), .Y(n3126) );
  MX2 U3451 ( .A(n3171), .B(n3172), .S0(n2699), .Y(n3170) );
  NOR2 U3452 ( .A(\uut/mult_mant/temp_product[12] ), .B(n3061), .Y(n3169) );
  OAI2BB2 U3453 ( .B0(n3173), .B1(n3066), .A0N(
        \uut/mult_mant/temp_product[11] ), .A1N(n3065), .Y(n3061) );
  NAND2B U3454 ( .AN(n2725), .B(n3128), .Y(n3066) );
  NOR2B U3455 ( .AN(n3174), .B(n2549), .Y(n3128) );
  MX2 U3456 ( .A(n3175), .B(n3176), .S0(n2699), .Y(n3174) );
  NOR2 U3457 ( .A(\uut/mult_mant/temp_product[11] ), .B(n3065), .Y(n3173) );
  OAI2BB2 U3458 ( .B0(n3177), .B1(n3070), .A0N(
        \uut/mult_mant/temp_product[10] ), .A1N(n3069), .Y(n3065) );
  NAND2B U3459 ( .AN(n2725), .B(n3130), .Y(n3070) );
  NOR2B U3460 ( .AN(n3178), .B(n2549), .Y(n3130) );
  MX2 U3461 ( .A(n3179), .B(n3180), .S0(n2699), .Y(n3178) );
  NOR2 U3462 ( .A(\uut/mult_mant/temp_product[10] ), .B(n3069), .Y(n3177) );
  OAI2BB2 U3463 ( .B0(n3181), .B1(n3074), .A0N(\uut/mult_mant/temp_product[9] ), .A1N(n3073), .Y(n3069) );
  NAND2B U3464 ( .AN(n2725), .B(n3132), .Y(n3074) );
  NOR2B U3465 ( .AN(n3182), .B(n2549), .Y(n3132) );
  MX2 U3466 ( .A(n3183), .B(n3184), .S0(n2699), .Y(n3182) );
  NOR2 U3467 ( .A(\uut/mult_mant/temp_product[9] ), .B(n3073), .Y(n3181) );
  OAI2BB2 U3468 ( .B0(n3185), .B1(n3078), .A0N(\uut/mult_mant/temp_product[8] ), .A1N(n3077), .Y(n3073) );
  NAND2B U3469 ( .AN(n2725), .B(n3134), .Y(n3078) );
  NOR2B U3470 ( .AN(n3186), .B(n2549), .Y(n3134) );
  MX2 U3471 ( .A(n3187), .B(n3188), .S0(n2699), .Y(n3186) );
  NOR2 U3472 ( .A(\uut/mult_mant/temp_product[8] ), .B(n3077), .Y(n3185) );
  OAI2BB2 U3473 ( .B0(n3189), .B1(n3082), .A0N(\uut/mult_mant/temp_product[7] ), .A1N(n3081), .Y(n3077) );
  NAND2 U3474 ( .A(n2643), .B(n3191), .Y(n3082) );
  NOR2 U3475 ( .A(\uut/mult_mant/temp_product[7] ), .B(n3081), .Y(n3189) );
  OAI2BB2 U3476 ( .B0(n3192), .B1(n3086), .A0N(\uut/mult_mant/temp_product[6] ), .A1N(n3085), .Y(n3081) );
  NAND2 U3477 ( .A(n3164), .B(n2643), .Y(n3086) );
  NOR2 U3478 ( .A(\uut/mult_mant/temp_product[6] ), .B(n3085), .Y(n3192) );
  OAI2BB2 U3479 ( .B0(n3193), .B1(n3090), .A0N(\uut/mult_mant/temp_product[5] ), .A1N(n3089), .Y(n3085) );
  NAND2 U3480 ( .A(n2643), .B(n3168), .Y(n3090) );
  NOR2 U3481 ( .A(\uut/mult_mant/temp_product[5] ), .B(n3089), .Y(n3193) );
  OAI2BB2 U3482 ( .B0(n3194), .B1(n3094), .A0N(\uut/mult_mant/temp_product[4] ), .A1N(n3093), .Y(n3089) );
  NAND2 U3483 ( .A(n3172), .B(n2643), .Y(n3094) );
  NOR2 U3484 ( .A(\uut/mult_mant/temp_product[4] ), .B(n3093), .Y(n3194) );
  OAI2BB2 U3485 ( .B0(n3097), .B1(n3195), .A0N(\uut/mult_mant/temp_product[3] ), .A1N(n3098), .Y(n3093) );
  NOR2 U3486 ( .A(n3098), .B(\uut/mult_mant/temp_product[3] ), .Y(n3195) );
  NOR2B U3487 ( .AN(n2643), .B(n3196), .Y(n3098) );
  INV U3488 ( .A(n3176), .Y(n3196) );
  AOI2BB2 U3489 ( .B0(\uut/mult_mant/temp_product[2] ), .B1(n3101), .A0N(n3197), .A1N(n3102), .Y(n3097) );
  NAND2 U3490 ( .A(n3180), .B(n2643), .Y(n3102) );
  NOR2 U3491 ( .A(\uut/mult_mant/temp_product[2] ), .B(n3101), .Y(n3197) );
  OAI2BB2 U3492 ( .B0(n3198), .B1(n3106), .A0N(n3105), .A1N(
        \uut/mult_mant/temp_product[1] ), .Y(n3101) );
  NAND2 U3493 ( .A(n3109), .B(\uut/mult_mant/temp_product[0] ), .Y(n3106) );
  NOR2B U3494 ( .AN(n3188), .B(n2642), .Y(n3109) );
  NOR2 U3495 ( .A(n3105), .B(\uut/mult_mant/temp_product[1] ), .Y(n3198) );
  NOR2B U3496 ( .AN(n2643), .B(n3199), .Y(n3105) );
  INV U3497 ( .A(n3184), .Y(n3199) );
  NOR2B U3498 ( .AN(n3200), .B(n2725), .Y(n3190) );
  AOI22 U3499 ( .A0(n3188), .A1(n2750), .B0(n3187), .B1(n2717), .Y(n3045) );
  AOI22 U3500 ( .A0(n3184), .A1(n2750), .B0(n3183), .B1(n2717), .Y(n3041) );
  AOI22 U3501 ( .A0(n3180), .A1(n2750), .B0(n3179), .B1(n2717), .Y(n3037) );
  AOI22 U3502 ( .A0(n2717), .A1(n3175), .B0(n2750), .B1(n3176), .Y(n3033) );
  AOI22 U3503 ( .A0(n3172), .A1(n2750), .B0(n3171), .B1(n2717), .Y(n3029) );
  AOI22 U3504 ( .A0(n2717), .A1(n3167), .B0(n2750), .B1(n3168), .Y(n3025) );
  AOI22 U3505 ( .A0(n3164), .A1(n2750), .B0(n3163), .B1(n2717), .Y(n3021) );
  AOI22 U3506 ( .A0(n2717), .A1(n3203), .B0(n2750), .B1(n3191), .Y(n3017) );
  NOR3B U3507 ( .AN(n2699), .B(n2725), .C(n2549), .Y(n3202) );
  AOI22 U3508 ( .A0(n2752), .A1(n3188), .B0(n3187), .B1(n2750), .Y(n3013) );
  AOI22 U3509 ( .A0(n2752), .A1(n3184), .B0(n3183), .B1(n2750), .Y(n3009) );
  AOI22 U3510 ( .A0(n2752), .A1(n3180), .B0(n3179), .B1(n2750), .Y(n3005) );
  AOI22 U3511 ( .A0(n2752), .A1(n3176), .B0(n2750), .B1(n3175), .Y(n3001) );
  AOI22 U3512 ( .A0(n2752), .A1(n3172), .B0(n3171), .B1(n2750), .Y(n2997) );
  AOI22 U3513 ( .A0(n2752), .A1(n3168), .B0(n2750), .B1(n3167), .Y(n2993) );
  AOI22 U3514 ( .A0(n2752), .A1(n3164), .B0(n3163), .B1(n2750), .Y(n2989) );
  AOI22 U3515 ( .A0(n2750), .A1(n3203), .B0(n2752), .B1(n3191), .Y(n2985) );
  NOR2B U3516 ( .AN(n3205), .B(n2699), .Y(n3201) );
  AOI22 U3517 ( .A0(n2645), .A1(n3188), .B0(n2752), .B1(n3187), .Y(n2981) );
  ADDF U3518 ( .A(n3207), .B(n3208), .CI(n3209), .S(n3187) );
  NOR2B U3519 ( .AN(\uut/mult_mant/in2_segment [0]), .B(n3210), .Y(n3188) );
  AOI22 U3520 ( .A0(n2645), .A1(n3184), .B0(n2752), .B1(n3183), .Y(n2977) );
  ADDF U3521 ( .A(n3211), .B(n3212), .CI(n3213), .S(n3183) );
  XOR2 U3522 ( .A(n3214), .B(n3215), .Y(n3184) );
  INV U3523 ( .A(n3216), .Y(n3215) );
  AOI22 U3524 ( .A0(n2645), .A1(n3180), .B0(n2752), .B1(n3179), .Y(n2973) );
  ADDF U3525 ( .A(n3217), .B(n3218), .CI(n3219), .S(n3179) );
  ADDF U3526 ( .A(n3220), .B(n3221), .CI(n3222), .S(n3180) );
  AOI22 U3527 ( .A0(n2645), .A1(n3176), .B0(n2752), .B1(n3175), .Y(n2969) );
  ADDF U3528 ( .A(n3223), .B(n3224), .CI(n3225), .S(n3175) );
  ADDF U3529 ( .A(n3226), .B(n3227), .CI(n3228), .S(n3176) );
  AOI22 U3530 ( .A0(n2645), .A1(n3172), .B0(n2752), .B1(n3171), .Y(n2965) );
  ADDF U3531 ( .A(n3229), .B(n3230), .CI(n3231), .S(n3171) );
  ADDF U3532 ( .A(n3232), .B(n3233), .CI(n3234), .S(n3172) );
  AOI22 U3533 ( .A0(n2645), .A1(n3168), .B0(n2752), .B1(n3167), .Y(n2961) );
  ADDF U3534 ( .A(n3235), .B(n3236), .CI(n3237), .S(n3167) );
  ADDF U3535 ( .A(n3238), .B(n3239), .CI(n3240), .S(n3168) );
  AOI22 U3536 ( .A0(n2645), .A1(n3164), .B0(n2752), .B1(n3163), .Y(n2957) );
  ADDF U3537 ( .A(n3241), .B(n3242), .CI(n3243), .S(n3163) );
  ADDF U3538 ( .A(n3244), .B(n3245), .CI(n3246), .S(n3164) );
  AOI22 U3539 ( .A0(n2752), .A1(n3203), .B0(n2645), .B1(n3191), .Y(n2953) );
  NOR2B U3540 ( .AN(n3200), .B(n2724), .Y(n3206) );
  NOR2B U3541 ( .AN(n3205), .B(n2698), .Y(n3204) );
  NOR2B U3542 ( .AN(n2549), .B(n2725), .Y(n3205) );
  NOR2 U3543 ( .A(n3160), .B(n2724), .Y(n3116) );
  AOI22 U3544 ( .A0(n3200), .A1(n3203), .B0(n3247), .B1(n3191), .Y(n3160) );
  ADDF U3545 ( .A(n3248), .B(n3249), .CI(n3250), .S(n3191) );
  NOR2B U3546 ( .AN(n2699), .B(n2549), .Y(n3247) );
  ADDF U3547 ( .A(n3241), .B(n3243), .CI(n3242), .CO(n3203) );
  ADDF U3548 ( .A(n3235), .B(n3236), .CI(n3237), .CO(n3242) );
  ADDF U3549 ( .A(n3251), .B(n3252), .CI(n3253), .S(n3237) );
  ADDF U3550 ( .A(n3254), .B(n3255), .CI(n3256), .CO(n3236) );
  ADDF U3551 ( .A(n3229), .B(n3231), .CI(n3230), .CO(n3235) );
  ADDF U3552 ( .A(n3257), .B(n3258), .CI(n3259), .CO(n3230) );
  ADDF U3553 ( .A(n3223), .B(n3224), .CI(n3225), .CO(n3231) );
  ADDF U3554 ( .A(n3257), .B(n3258), .CI(n3259), .S(n3225) );
  ADDF U3555 ( .A(n3260), .B(n3261), .CI(n3262), .S(n3259) );
  ADDF U3556 ( .A(n3263), .B(n3264), .CI(n3265), .CO(n3258) );
  ADDF U3557 ( .A(n3266), .B(n3267), .CI(n3268), .CO(n3257) );
  ADDF U3558 ( .A(n3269), .B(n3270), .CI(n3271), .CO(n3224) );
  ADDF U3559 ( .A(n3217), .B(n3219), .CI(n3218), .CO(n3223) );
  ADDF U3560 ( .A(n3211), .B(n3213), .CI(n3212), .CO(n3218) );
  ADDF U3561 ( .A(n3207), .B(n3209), .CI(n3208), .CO(n3212) );
  ADDF U3562 ( .A(n3248), .B(n3249), .CI(n3250), .CO(n3208) );
  ADDF U3563 ( .A(n3272), .B(n3273), .CI(n3274), .S(n3250) );
  ADDF U3564 ( .A(n3275), .B(n3276), .CI(n3277), .CO(n3249) );
  ADDF U3565 ( .A(n3244), .B(n3246), .CI(n3245), .CO(n3248) );
  ADDF U3566 ( .A(n3238), .B(n3239), .CI(n3240), .CO(n3245) );
  ADDF U3567 ( .A(n3278), .B(n3279), .CI(n3280), .S(n3240) );
  ADDF U3568 ( .A(n3281), .B(n3282), .CI(n3283), .CO(n3239) );
  ADDF U3569 ( .A(n3232), .B(n3234), .CI(n3233), .CO(n3238) );
  ADDF U3570 ( .A(n3226), .B(n3227), .CI(n3228), .CO(n3233) );
  ADDF U3571 ( .A(n3220), .B(n3221), .CI(n3222), .CO(n3228) );
  NOR2B U3572 ( .AN(\uut/mult_mant/in2_segment [2]), .B(n3210), .Y(n3222) );
  XOR2 U3573 ( .A(n3284), .B(n3285), .Y(n3221) );
  INV U3574 ( .A(n3286), .Y(n3285) );
  NOR2B U3575 ( .AN(n3214), .B(n3216), .Y(n3220) );
  NAND2 U3576 ( .A(\uut/mult_mant/in2_segment [1]), .B(
        \uut/mult_mant/in1_segment [0]), .Y(n3216) );
  NOR2B U3577 ( .AN(\uut/mult_mant/in1_segment [1]), .B(n3287), .Y(n3214) );
  INV U3578 ( .A(\uut/mult_mant/in2_segment [0]), .Y(n3287) );
  XOR2 U3579 ( .A(n3288), .B(n3289), .Y(n3227) );
  INV U3580 ( .A(n3290), .Y(n3289) );
  ADDF U3581 ( .A(n3291), .B(n3292), .CI(n3293), .S(n3226) );
  ADDF U3582 ( .A(n3291), .B(n3292), .CI(n3293), .CO(n3234) );
  NOR2B U3583 ( .AN(\uut/mult_mant/in2_segment [3]), .B(n3210), .Y(n3293) );
  INV U3584 ( .A(\uut/mult_mant/in1_segment [0]), .Y(n3210) );
  NOR2B U3585 ( .AN(\uut/mult_mant/in1_segment [1]), .B(n3294), .Y(n3292) );
  NOR2B U3586 ( .AN(n3284), .B(n3286), .Y(n3291) );
  NAND2 U3587 ( .A(\uut/mult_mant/in1_segment [2]), .B(
        \uut/mult_mant/in2_segment [0]), .Y(n3286) );
  NOR2B U3588 ( .AN(\uut/mult_mant/in1_segment [1]), .B(n3295), .Y(n3284) );
  INV U3589 ( .A(\uut/mult_mant/in2_segment [1]), .Y(n3295) );
  ADDF U3590 ( .A(n3281), .B(n3282), .CI(n3283), .S(n3232) );
  XOR2 U3591 ( .A(n3296), .B(n3297), .Y(n3283) );
  INV U3592 ( .A(n3298), .Y(n3297) );
  NOR2B U3593 ( .AN(n3288), .B(n3290), .Y(n3282) );
  NAND2 U3594 ( .A(\uut/mult_mant/in2_segment [0]), .B(
        \uut/mult_mant/in1_segment [3]), .Y(n3290) );
  NOR2B U3595 ( .AN(\uut/mult_mant/in2_segment [1]), .B(n3299), .Y(n3288) );
  INV U3596 ( .A(\uut/mult_mant/in1_segment [2]), .Y(n3299) );
  ADDF U3597 ( .A(n3300), .B(n3301), .CI(n3302), .S(n3281) );
  ADDF U3598 ( .A(n3278), .B(n3279), .CI(n3280), .CO(n3246) );
  ADDF U3599 ( .A(n3303), .B(n3304), .CI(n3305), .S(n3280) );
  XOR2 U3600 ( .A(n3306), .B(n3307), .Y(n3279) );
  INV U3601 ( .A(n3308), .Y(n3307) );
  ADDF U3602 ( .A(n3309), .B(n3310), .CI(n3311), .S(n3278) );
  ADDF U3603 ( .A(n3275), .B(n3276), .CI(n3277), .S(n3244) );
  ADDF U3604 ( .A(n3312), .B(n3313), .CI(n3314), .S(n3277) );
  ADDF U3605 ( .A(n3303), .B(n3304), .CI(n3305), .CO(n3276) );
  ADDF U3606 ( .A(n3300), .B(n3301), .CI(n3302), .CO(n3305) );
  NOR2B U3607 ( .AN(\uut/mult_mant/in1_segment [2]), .B(n3294), .Y(n3302) );
  INV U3608 ( .A(\uut/mult_mant/in2_segment [2]), .Y(n3294) );
  NOR2B U3609 ( .AN(\uut/mult_mant/in1_segment [1]), .B(n3315), .Y(n3301) );
  NOR2B U3610 ( .AN(\uut/mult_mant/in1_segment [0]), .B(n3316), .Y(n3300) );
  NOR2B U3611 ( .AN(\uut/mult_mant/in1_segment [0]), .B(n3317), .Y(n3304) );
  NOR2B U3612 ( .AN(n3296), .B(n3298), .Y(n3303) );
  NAND2 U3613 ( .A(\uut/mult_mant/in2_segment [0]), .B(
        \uut/mult_mant/in1_segment [4]), .Y(n3298) );
  NOR2B U3614 ( .AN(\uut/mult_mant/in2_segment [1]), .B(n3318), .Y(n3296) );
  ADDF U3615 ( .A(n3319), .B(n3320), .CI(n3321), .S(n3275) );
  ADDF U3616 ( .A(n3272), .B(n3273), .CI(n3274), .CO(n3209) );
  ADDF U3617 ( .A(n3322), .B(n3323), .CI(n3324), .S(n3274) );
  ADDF U3618 ( .A(n3325), .B(n3326), .CI(n3327), .S(n3273) );
  ADDF U3619 ( .A(n3312), .B(n3313), .CI(n3314), .CO(n3272) );
  ADDF U3620 ( .A(n3309), .B(n3310), .CI(n3311), .CO(n3314) );
  NOR2B U3621 ( .AN(\uut/mult_mant/in1_segment [1]), .B(n3316), .Y(n3311) );
  NOR2B U3622 ( .AN(\uut/mult_mant/in2_segment [2]), .B(n3318), .Y(n3310) );
  NOR2B U3623 ( .AN(\uut/mult_mant/in1_segment [2]), .B(n3315), .Y(n3309) );
  INV U3624 ( .A(\uut/mult_mant/in2_segment [3]), .Y(n3315) );
  ADDF U3625 ( .A(n3328), .B(n3329), .CI(n3330), .S(n3313) );
  XOR2 U3626 ( .A(n3331), .B(n3332), .Y(n3312) );
  INV U3627 ( .A(n3333), .Y(n3332) );
  ADDF U3628 ( .A(n3334), .B(n3335), .CI(n3336), .S(n3207) );
  ADDF U3629 ( .A(n3334), .B(n3336), .CI(n3335), .CO(n3213) );
  ADDF U3630 ( .A(n3325), .B(n3326), .CI(n3327), .CO(n3335) );
  ADDF U3631 ( .A(n3319), .B(n3320), .CI(n3321), .CO(n3327) );
  NOR2B U3632 ( .AN(\uut/mult_mant/in1_segment [1]), .B(n3317), .Y(n3321) );
  NOR2B U3633 ( .AN(\uut/mult_mant/in1_segment [0]), .B(n3337), .Y(n3320) );
  NOR2B U3634 ( .AN(n3306), .B(n3308), .Y(n3319) );
  NAND2 U3635 ( .A(\uut/mult_mant/in2_segment [0]), .B(
        \uut/mult_mant/in1_segment [5]), .Y(n3308) );
  NOR2B U3636 ( .AN(\uut/mult_mant/in2_segment [1]), .B(n3338), .Y(n3306) );
  ADDF U3637 ( .A(n3339), .B(n3340), .CI(n3341), .S(n3326) );
  XOR2 U3638 ( .A(n3342), .B(n3343), .Y(n3325) );
  INV U3639 ( .A(n3344), .Y(n3343) );
  ADDF U3640 ( .A(n3345), .B(n3346), .CI(n3347), .S(n3336) );
  ADDF U3641 ( .A(n3348), .B(n3349), .CI(n3350), .S(n3334) );
  ADDF U3642 ( .A(n3351), .B(n3352), .CI(n3353), .S(n3211) );
  ADDF U3643 ( .A(n3351), .B(n3352), .CI(n3353), .CO(n3219) );
  ADDF U3644 ( .A(n3354), .B(n3355), .CI(n3356), .S(n3353) );
  ADDF U3645 ( .A(n3345), .B(n3346), .CI(n3347), .CO(n3352) );
  ADDF U3646 ( .A(n3322), .B(n3323), .CI(n3324), .CO(n3347) );
  ADDF U3647 ( .A(n3328), .B(n3329), .CI(n3330), .CO(n3324) );
  NOR2B U3648 ( .AN(\uut/mult_mant/in1_segment [2]), .B(n3316), .Y(n3330) );
  NOR2B U3649 ( .AN(\uut/mult_mant/in2_segment [3]), .B(n3318), .Y(n3329) );
  INV U3650 ( .A(\uut/mult_mant/in1_segment [3]), .Y(n3318) );
  NOR2B U3651 ( .AN(\uut/mult_mant/in2_segment [2]), .B(n3338), .Y(n3328) );
  ADDF U3652 ( .A(n3357), .B(n3358), .CI(n3359), .S(n3323) );
  NOR2B U3653 ( .AN(n3331), .B(n3333), .Y(n3322) );
  NAND2 U3654 ( .A(\uut/mult_mant/in2_segment [0]), .B(
        \uut/mult_mant/in1_segment [6]), .Y(n3333) );
  NOR2B U3655 ( .AN(\uut/mult_mant/in2_segment [1]), .B(n3360), .Y(n3331) );
  XOR2 U3656 ( .A(n3361), .B(n3362), .Y(n3346) );
  INV U3657 ( .A(n3363), .Y(n3362) );
  ADDF U3658 ( .A(n3364), .B(n3365), .CI(n3366), .S(n3345) );
  ADDF U3659 ( .A(n3367), .B(n3368), .CI(n3369), .S(n3351) );
  ADDF U3660 ( .A(n3269), .B(n3270), .CI(n3271), .S(n3217) );
  ADDF U3661 ( .A(n3354), .B(n3355), .CI(n3356), .CO(n3271) );
  ADDF U3662 ( .A(n3370), .B(n3371), .CI(n3372), .CO(n3356) );
  ADDF U3663 ( .A(n3373), .B(n3374), .CI(n3375), .S(n3355) );
  NOR2B U3664 ( .AN(n3361), .B(n3363), .Y(n3354) );
  NAND2 U3665 ( .A(\uut/mult_mant/in2_segment [2]), .B(
        \uut/mult_mant/in1_segment [6]), .Y(n3363) );
  NOR2B U3666 ( .AN(\uut/mult_mant/in2_segment [1]), .B(n3376), .Y(n3361) );
  ADDF U3667 ( .A(n3367), .B(n3369), .CI(n3368), .CO(n3270) );
  ADDF U3668 ( .A(n3348), .B(n3349), .CI(n3350), .CO(n3368) );
  ADDF U3669 ( .A(n3357), .B(n3358), .CI(n3359), .CO(n3350) );
  NOR2B U3670 ( .AN(\uut/mult_mant/in2_segment [3]), .B(n3338), .Y(n3359) );
  NOR2B U3671 ( .AN(\uut/mult_mant/in1_segment [3]), .B(n3316), .Y(n3358) );
  INV U3672 ( .A(\uut/mult_mant/in2_segment [4]), .Y(n3316) );
  NOR2B U3673 ( .AN(\uut/mult_mant/in2_segment [2]), .B(n3360), .Y(n3357) );
  ADDF U3674 ( .A(n3339), .B(n3340), .CI(n3341), .CO(n3349) );
  NOR2B U3675 ( .AN(\uut/mult_mant/in1_segment [0]), .B(n3377), .Y(n3341) );
  NOR2B U3676 ( .AN(\uut/mult_mant/in1_segment [1]), .B(n3337), .Y(n3340) );
  NOR2B U3677 ( .AN(\uut/mult_mant/in1_segment [2]), .B(n3317), .Y(n3339) );
  ADDF U3678 ( .A(n3370), .B(n3371), .CI(n3372), .S(n3348) );
  NOR2B U3679 ( .AN(\uut/mult_mant/in2_segment [4]), .B(n3338), .Y(n3372) );
  INV U3680 ( .A(\uut/mult_mant/in1_segment [4]), .Y(n3338) );
  NOR2B U3681 ( .AN(\uut/mult_mant/in1_segment [2]), .B(n3337), .Y(n3371) );
  NOR2B U3682 ( .AN(\uut/mult_mant/in2_segment [3]), .B(n3360), .Y(n3370) );
  ADDF U3683 ( .A(n3364), .B(n3365), .CI(n3366), .CO(n3369) );
  NOR2B U3684 ( .AN(\uut/mult_mant/in1_segment [3]), .B(n3317), .Y(n3366) );
  NOR2B U3685 ( .AN(\uut/mult_mant/in1_segment [1]), .B(n3377), .Y(n3365) );
  NOR2B U3686 ( .AN(n3342), .B(n3344), .Y(n3364) );
  NAND2 U3687 ( .A(\uut/mult_mant/in2_segment [0]), .B(
        \uut/mult_mant/in1_segment [7]), .Y(n3344) );
  NOR2B U3688 ( .AN(\uut/mult_mant/in2_segment [1]), .B(n3378), .Y(n3342) );
  ADDF U3689 ( .A(n3379), .B(n3380), .CI(n3381), .S(n3367) );
  ADDF U3690 ( .A(n3266), .B(n3268), .CI(n3267), .S(n3269) );
  ADDF U3691 ( .A(n3379), .B(n3380), .CI(n3381), .CO(n3267) );
  NOR2B U3692 ( .AN(\uut/mult_mant/in1_segment [2]), .B(n3377), .Y(n3381) );
  NOR2B U3693 ( .AN(\uut/mult_mant/in1_segment [3]), .B(n3337), .Y(n3380) );
  NOR2B U3694 ( .AN(\uut/mult_mant/in1_segment [4]), .B(n3317), .Y(n3379) );
  INV U3695 ( .A(\uut/mult_mant/in2_segment [5]), .Y(n3317) );
  ADDF U3696 ( .A(n3263), .B(n3264), .CI(n3265), .S(n3268) );
  ADDF U3697 ( .A(n3373), .B(n3374), .CI(n3375), .CO(n3265) );
  NOR2B U3698 ( .AN(\uut/mult_mant/in2_segment [2]), .B(n3376), .Y(n3375) );
  NOR2B U3699 ( .AN(\uut/mult_mant/in2_segment [4]), .B(n3360), .Y(n3374) );
  NOR2B U3700 ( .AN(\uut/mult_mant/in2_segment [3]), .B(n3378), .Y(n3373) );
  NOR2B U3701 ( .AN(\uut/mult_mant/in1_segment [3]), .B(n3377), .Y(n3264) );
  NOR2B U3702 ( .AN(\uut/mult_mant/in2_segment [5]), .B(n3360), .Y(n3263) );
  INV U3703 ( .A(\uut/mult_mant/in1_segment [5]), .Y(n3360) );
  ADDF U3704 ( .A(n3382), .B(n3383), .CI(n3384), .S(n3266) );
  ADDF U3705 ( .A(n3254), .B(n3256), .CI(n3255), .S(n3229) );
  ADDF U3706 ( .A(n3385), .B(n3386), .CI(n3387), .CO(n3255) );
  ADDF U3707 ( .A(n3260), .B(n3261), .CI(n3262), .CO(n3256) );
  ADDF U3708 ( .A(n3382), .B(n3383), .CI(n3384), .CO(n3262) );
  NOR2B U3709 ( .AN(\uut/mult_mant/in2_segment [3]), .B(n3376), .Y(n3384) );
  NOR2B U3710 ( .AN(\uut/mult_mant/in1_segment [4]), .B(n3337), .Y(n3383) );
  NOR2B U3711 ( .AN(\uut/mult_mant/in2_segment [4]), .B(n3378), .Y(n3382) );
  NOR2B U3712 ( .AN(\uut/mult_mant/in1_segment [4]), .B(n3377), .Y(n3261) );
  ADDF U3713 ( .A(n3385), .B(n3386), .CI(n3387), .S(n3260) );
  NOR2B U3714 ( .AN(\uut/mult_mant/in1_segment [5]), .B(n3337), .Y(n3387) );
  INV U3715 ( .A(\uut/mult_mant/in2_segment [6]), .Y(n3337) );
  NOR2B U3716 ( .AN(\uut/mult_mant/in2_segment [4]), .B(n3376), .Y(n3386) );
  NOR2B U3717 ( .AN(\uut/mult_mant/in2_segment [5]), .B(n3378), .Y(n3385) );
  ADDF U3718 ( .A(n3388), .B(n3389), .CI(n3390), .S(n3254) );
  ADDF U3719 ( .A(n3251), .B(n3252), .CI(n3253), .CO(n3243) );
  ADDF U3720 ( .A(n3388), .B(n3389), .CI(n3390), .CO(n3253) );
  NOR2B U3721 ( .AN(\uut/mult_mant/in1_segment [5]), .B(n3377), .Y(n3390) );
  NOR2B U3722 ( .AN(\uut/mult_mant/in2_segment [5]), .B(n3376), .Y(n3389) );
  NOR2B U3723 ( .AN(\uut/mult_mant/in2_segment [6]), .B(n3378), .Y(n3388) );
  INV U3724 ( .A(\uut/mult_mant/in1_segment [6]), .Y(n3378) );
  NOR2B U3725 ( .AN(\uut/mult_mant/in1_segment [6]), .B(n3377), .Y(n3252) );
  NOR2B U3726 ( .AN(\uut/mult_mant/in2_segment [6]), .B(n3376), .Y(n3251) );
  INV U3727 ( .A(\uut/mult_mant/in1_segment [7]), .Y(n3376) );
  NOR2B U3728 ( .AN(\uut/mult_mant/in1_segment [7]), .B(n3377), .Y(n3241) );
  INV U3729 ( .A(\uut/mult_mant/in2_segment [7]), .Y(n3377) );
  NOR2 U3730 ( .A(n2549), .B(n2699), .Y(n3200) );
  NOR2 U3731 ( .A(n3391), .B(n3392), .Y(n3112) );
  INV U3732 ( .A(\uut/mult_mant/temp_product[47] ), .Y(n3111) );
  NOR2B U3733 ( .AN(in1_row[3]), .B(n3393), .Y(n4962) );
  NOR2B U3734 ( .AN(in1_row[2]), .B(n3393), .Y(n4963) );
  NOR2B U3735 ( .AN(in1_row[1]), .B(n3393), .Y(n4964) );
  NOR2B U3736 ( .AN(in1_row[0]), .B(n3393), .Y(n4965) );
  OR4 U3737 ( .A(in1_row_q[3]), .B(in1_row_q[2]), .C(in1_row_q[1]), .D(
        in1_row_q[0]), .Y(n3393) );
  NOR2B U3738 ( .AN(in1_col[3]), .B(n3394), .Y(n4966) );
  NOR2B U3739 ( .AN(in1_col[2]), .B(n3394), .Y(n4967) );
  NOR2B U3740 ( .AN(in1_col[1]), .B(n3394), .Y(n4968) );
  NOR2B U3741 ( .AN(in1_col[0]), .B(n3394), .Y(n4969) );
  OR4 U3742 ( .A(in1_col_q[3]), .B(in1_col_q[2]), .C(in1_col_q[1]), .D(
        in1_col_q[0]), .Y(n3394) );
  NOR2B U3743 ( .AN(in2_row[3]), .B(n3395), .Y(n4970) );
  NOR2B U3744 ( .AN(in2_row[2]), .B(n3395), .Y(n4971) );
  NOR2B U3745 ( .AN(in2_row[1]), .B(n3395), .Y(n4972) );
  NOR2B U3746 ( .AN(in2_row[0]), .B(n3395), .Y(n4973) );
  OR4 U3747 ( .A(in2_row_q[3]), .B(in2_row_q[2]), .C(in2_row_q[1]), .D(
        in2_row_q[0]), .Y(n3395) );
  NOR2B U3748 ( .AN(in2_col[3]), .B(n3396), .Y(n4974) );
  NOR2B U3749 ( .AN(in2_col[2]), .B(n3396), .Y(n4975) );
  NOR2B U3750 ( .AN(in2_col[1]), .B(n3396), .Y(n4976) );
  NOR2B U3751 ( .AN(in2_col[0]), .B(n3396), .Y(n4977) );
  OR4 U3752 ( .A(in2_col_q[3]), .B(in2_col_q[2]), .C(in2_col_q[1]), .D(
        in2_col_q[0]), .Y(n3396) );
  NAND4 U3753 ( .A(n3397), .B(n3398), .C(n3399), .D(n3400), .Y(out_seg[0]) );
  AOI22 U3754 ( .A0(out_sel[6]), .A1(bit6[0]), .B0(out_sel[5]), .B1(bit5[0]), 
        .Y(n3400) );
  AOI22 U3755 ( .A0(out_sel[4]), .A1(bit4[0]), .B0(out_sel[3]), .B1(bit3[0]), 
        .Y(n3399) );
  AOI22 U3756 ( .A0(out_sel[2]), .A1(bit2[0]), .B0(out_sel[1]), .B1(bit1[0]), 
        .Y(n3398) );
  AOI22 U3757 ( .A0(out_sel[7]), .A1(bit7[0]), .B0(out_sel[0]), .B1(bit0[0]), 
        .Y(n3397) );
  NAND4 U3758 ( .A(n3401), .B(n3402), .C(n3403), .D(n3404), .Y(out_seg[1]) );
  AOI22 U3759 ( .A0(out_sel[6]), .A1(bit6[1]), .B0(out_sel[5]), .B1(bit5[1]), 
        .Y(n3404) );
  AOI22 U3760 ( .A0(out_sel[4]), .A1(bit4[1]), .B0(out_sel[3]), .B1(bit3[1]), 
        .Y(n3403) );
  AOI22 U3761 ( .A0(out_sel[2]), .A1(bit2[1]), .B0(out_sel[1]), .B1(bit1[1]), 
        .Y(n3402) );
  AOI22 U3762 ( .A0(out_sel[7]), .A1(bit7[1]), .B0(out_sel[0]), .B1(bit0[1]), 
        .Y(n3401) );
  NAND4 U3763 ( .A(n3405), .B(n3406), .C(n3407), .D(n3408), .Y(out_seg[2]) );
  AOI22 U3764 ( .A0(out_sel[6]), .A1(bit6[2]), .B0(out_sel[5]), .B1(bit5[2]), 
        .Y(n3408) );
  AOI22 U3765 ( .A0(out_sel[4]), .A1(bit4[2]), .B0(out_sel[3]), .B1(bit3[2]), 
        .Y(n3407) );
  AOI22 U3766 ( .A0(out_sel[2]), .A1(bit2[2]), .B0(out_sel[1]), .B1(bit1[2]), 
        .Y(n3406) );
  AOI22 U3767 ( .A0(out_sel[7]), .A1(bit7[2]), .B0(out_sel[0]), .B1(bit0[2]), 
        .Y(n3405) );
  NAND4 U3768 ( .A(n3409), .B(n3410), .C(n3411), .D(n3412), .Y(out_seg[3]) );
  AOI22 U3769 ( .A0(out_sel[6]), .A1(bit6[3]), .B0(out_sel[5]), .B1(bit5[3]), 
        .Y(n3412) );
  AOI22 U3770 ( .A0(out_sel[4]), .A1(bit4[3]), .B0(out_sel[3]), .B1(bit3[3]), 
        .Y(n3411) );
  AOI22 U3771 ( .A0(out_sel[2]), .A1(bit2[3]), .B0(out_sel[1]), .B1(bit1[3]), 
        .Y(n3410) );
  AOI22 U3772 ( .A0(out_sel[7]), .A1(bit7[3]), .B0(out_sel[0]), .B1(bit0[3]), 
        .Y(n3409) );
  NAND4 U3773 ( .A(n3413), .B(n3414), .C(n3415), .D(n3416), .Y(out_seg[4]) );
  AOI22 U3774 ( .A0(out_sel[6]), .A1(bit6[4]), .B0(out_sel[5]), .B1(bit5[4]), 
        .Y(n3416) );
  AOI22 U3775 ( .A0(out_sel[4]), .A1(bit4[4]), .B0(out_sel[3]), .B1(bit3[4]), 
        .Y(n3415) );
  AOI22 U3776 ( .A0(out_sel[2]), .A1(bit2[4]), .B0(out_sel[1]), .B1(bit1[4]), 
        .Y(n3414) );
  AOI22 U3777 ( .A0(out_sel[7]), .A1(bit7[4]), .B0(out_sel[0]), .B1(bit0[4]), 
        .Y(n3413) );
  NAND4 U3778 ( .A(n3417), .B(n3418), .C(n3419), .D(n3420), .Y(out_seg[5]) );
  AOI22 U3779 ( .A0(out_sel[6]), .A1(bit6[5]), .B0(out_sel[5]), .B1(bit5[5]), 
        .Y(n3420) );
  AOI22 U3780 ( .A0(out_sel[4]), .A1(bit4[5]), .B0(out_sel[3]), .B1(bit3[5]), 
        .Y(n3419) );
  AOI22 U3781 ( .A0(out_sel[2]), .A1(bit2[5]), .B0(out_sel[1]), .B1(bit1[5]), 
        .Y(n3418) );
  AOI22 U3782 ( .A0(out_sel[7]), .A1(bit7[5]), .B0(out_sel[0]), .B1(bit0[5]), 
        .Y(n3417) );
  NAND4 U3783 ( .A(n3421), .B(n3422), .C(n3423), .D(n3424), .Y(out_seg[6]) );
  AOI22 U3784 ( .A0(out_sel[6]), .A1(bit6[6]), .B0(out_sel[5]), .B1(bit5[6]), 
        .Y(n3424) );
  NOR2B U3785 ( .AN(n3425), .B(n3426), .Y(n5002) );
  NOR3B U3786 ( .AN(out_sel_cnt[2]), .B(out_sel_cnt[0]), .C(n3427), .Y(n5001)
         );
  AOI22 U3787 ( .A0(out_sel[4]), .A1(bit4[6]), .B0(out_sel[3]), .B1(bit3[6]), 
        .Y(n3423) );
  NOR2B U3788 ( .AN(n3428), .B(n3426), .Y(n5004) );
  NOR2B U3789 ( .AN(n3425), .B(out_sel_cnt[0]), .Y(n5003) );
  NOR2B U3790 ( .AN(out_sel_cnt[2]), .B(out_sel_cnt[1]), .Y(n3425) );
  AOI22 U3791 ( .A0(out_sel[2]), .A1(bit2[6]), .B0(out_sel[1]), .B1(bit1[6]), 
        .Y(n3422) );
  NOR2B U3792 ( .AN(n3429), .B(n3426), .Y(n5006) );
  NOR2B U3793 ( .AN(n3428), .B(out_sel_cnt[0]), .Y(n5005) );
  NOR2 U3794 ( .A(out_sel_cnt[2]), .B(n3427), .Y(n3428) );
  AOI22 U3795 ( .A0(out_sel[7]), .A1(bit7[6]), .B0(out_sel[0]), .B1(bit0[6]), 
        .Y(n3421) );
  NOR3B U3796 ( .AN(out_sel_cnt[2]), .B(n3427), .C(n3426), .Y(n4987) );
  INV U3797 ( .A(out_sel_cnt[0]), .Y(n3426) );
  INV U3798 ( .A(out_sel_cnt[1]), .Y(n3427) );
  NOR2 U3799 ( .A(enter), .B(n3430), .Y(n2497) );
  XNOR2 U3800 ( .A(input1_cnt[0]), .B(n2771), .Y(n3430) );
  NOR2 U3801 ( .A(enter), .B(n3431), .Y(n2495) );
  XNOR2 U3802 ( .A(input1_cnt[1]), .B(n3432), .Y(n3431) );
  NOR2 U3803 ( .A(enter), .B(n3433), .Y(n2494) );
  XNOR2 U3804 ( .A(input1_cnt[2]), .B(n3434), .Y(n3433) );
  NOR2B U3805 ( .AN(n3432), .B(n3435), .Y(n3434) );
  INV U3806 ( .A(input1_cnt[1]), .Y(n3435) );
  NOR2 U3807 ( .A(n2772), .B(n3437), .Y(n3432) );
  NOR2 U3808 ( .A(enter), .B(n3438), .Y(n2493) );
  AOI21 U3809 ( .A0(n2771), .A1(n2561), .B0(input1_cnt[3]), .Y(n3438) );
  NOR2 U3810 ( .A(enter), .B(n3440), .Y(n2491) );
  XNOR2 U3811 ( .A(input2_cnt[0]), .B(n2769), .Y(n3440) );
  NOR2 U3812 ( .A(enter), .B(n3441), .Y(n2489) );
  XNOR2 U3813 ( .A(input2_cnt[1]), .B(n3442), .Y(n3441) );
  NOR2 U3814 ( .A(enter), .B(n3443), .Y(n2488) );
  XNOR2 U3815 ( .A(input2_cnt[2]), .B(n3444), .Y(n3443) );
  NOR2B U3816 ( .AN(n3442), .B(n3445), .Y(n3444) );
  INV U3817 ( .A(input2_cnt[1]), .Y(n3445) );
  NOR2 U3818 ( .A(n2770), .B(n3447), .Y(n3442) );
  NOR2 U3819 ( .A(enter), .B(n3448), .Y(n2487) );
  AOI21 U3820 ( .A0(n2769), .A1(n2559), .B0(input2_cnt[3]), .Y(n3448) );
  NAND2B U3821 ( .AN(n3450), .B(n2762), .Y(n2485) );
  MX2 U3822 ( .A(\uut/mult_ready ), .B(n2767), .S0(n2787), .Y(n3450) );
  OAI2BB2 U3823 ( .B0(n3451), .B1(n3452), .A0N(n2790), .A1N(n3453), .Y(n2484)
         );
  NOR2 U3824 ( .A(n2791), .B(n3454), .Y(n3451) );
  NOR2B U3825 ( .AN(n2697), .B(n2541), .Y(n3454) );
  MX2 U3826 ( .A(n3455), .B(n3456), .S0(\uut/mult_mant/mult8_cnt[2] ), .Y(
        n2483) );
  OAI21 U3827 ( .A0(n3457), .A1(n3458), .B0(n3459), .Y(n2482) );
  NOR2 U3828 ( .A(n2697), .B(n3456), .Y(n3457) );
  OAI21 U3829 ( .A0(n3460), .A1(n2696), .B0(n3461), .Y(n3456) );
  OAI211 U3830 ( .A0(n2698), .A1(n3461), .B0(n3459), .C0(n3462), .Y(n2481) );
  OAI211 U3831 ( .A0(n3463), .A1(n3464), .B0(n2790), .C0(n3458), .Y(n3462) );
  NOR2 U3832 ( .A(n2541), .B(n3452), .Y(n3464) );
  NOR2B U3833 ( .AN(n3453), .B(\uut/mult_mant/mult8_cnt[2] ), .Y(n3463) );
  NAND2 U3834 ( .A(n3455), .B(n3465), .Y(n3459) );
  OAI222 U3835 ( .A0(n3466), .A1(n3467), .B0(n2548), .B1(n3461), .C0(n3468), 
        .C1(n3469), .Y(n2480) );
  INV U3836 ( .A(n3455), .Y(n3468) );
  NOR2B U3837 ( .AN(n3460), .B(n3467), .Y(n3455) );
  INV U3838 ( .A(n2790), .Y(n3467) );
  OAI2BB2 U3839 ( .B0(n3461), .B1(n2724), .A0N(n2790), .A1N(n3470), .Y(n2479)
         );
  NOR2B U3840 ( .AN(n2697), .B(n2791), .Y(n2790) );
  INV U3841 ( .A(n2791), .Y(n3461) );
  NOR2 U3842 ( .A(n2787), .B(n2783), .Y(n2791) );
  MX2 U3843 ( .A(\uut/mult_mant/in1_segment [0]), .B(n3472), .S0(n2783), .Y(
        n2478) );
  INV U3844 ( .A(n3473), .Y(n3472) );
  AOI222 U3845 ( .A0(n2655), .A1(\uut/mult_mant/c1 [0]), .B0(n2653), .B1(
        \uut/mult_mant/b1 [0]), .C0(n2661), .C1(\uut/mult_mant/a1 [0]), .Y(
        n3473) );
  MX2 U3846 ( .A(\uut/mult_mant/in1_segment [1]), .B(n3477), .S0(n2783), .Y(
        n2477) );
  INV U3847 ( .A(n3478), .Y(n3477) );
  AOI222 U3848 ( .A0(n2655), .A1(\uut/mult_mant/c1 [1]), .B0(n2653), .B1(
        \uut/mult_mant/b1 [1]), .C0(n2661), .C1(\uut/mult_mant/a1 [1]), .Y(
        n3478) );
  MX2 U3849 ( .A(\uut/mult_mant/in1_segment [2]), .B(n3479), .S0(n2783), .Y(
        n2476) );
  INV U3850 ( .A(n3480), .Y(n3479) );
  AOI222 U3851 ( .A0(n2655), .A1(\uut/mult_mant/c1 [2]), .B0(n2653), .B1(
        \uut/mult_mant/b1 [2]), .C0(n2661), .C1(\uut/mult_mant/a1 [2]), .Y(
        n3480) );
  MX2 U3852 ( .A(\uut/mult_mant/in1_segment [3]), .B(n3481), .S0(n2783), .Y(
        n2475) );
  INV U3853 ( .A(n3482), .Y(n3481) );
  AOI222 U3854 ( .A0(n2655), .A1(\uut/mult_mant/c1 [3]), .B0(n2653), .B1(
        \uut/mult_mant/b1 [3]), .C0(n2661), .C1(\uut/mult_mant/a1 [3]), .Y(
        n3482) );
  MX2 U3855 ( .A(\uut/mult_mant/in1_segment [4]), .B(n3483), .S0(n2783), .Y(
        n2474) );
  INV U3856 ( .A(n3484), .Y(n3483) );
  AOI222 U3857 ( .A0(n2655), .A1(\uut/mult_mant/c1 [4]), .B0(n2653), .B1(
        \uut/mult_mant/b1 [4]), .C0(n2661), .C1(\uut/mult_mant/a1 [4]), .Y(
        n3484) );
  MX2 U3858 ( .A(\uut/mult_mant/in1_segment [5]), .B(n3485), .S0(n2783), .Y(
        n2473) );
  INV U3859 ( .A(n3486), .Y(n3485) );
  AOI222 U3860 ( .A0(n2655), .A1(\uut/mult_mant/c1 [5]), .B0(n2653), .B1(
        \uut/mult_mant/b1 [5]), .C0(n2661), .C1(\uut/mult_mant/a1 [5]), .Y(
        n3486) );
  MX2 U3861 ( .A(\uut/mult_mant/in1_segment [6]), .B(n3487), .S0(n2783), .Y(
        n2472) );
  INV U3862 ( .A(n3488), .Y(n3487) );
  AOI222 U3863 ( .A0(n2655), .A1(\uut/mult_mant/c1 [6]), .B0(n2653), .B1(
        \uut/mult_mant/b1 [6]), .C0(n2661), .C1(\uut/mult_mant/a1 [6]), .Y(
        n3488) );
  MX2 U3864 ( .A(\uut/mult_mant/in1_segment [7]), .B(n3489), .S0(n2783), .Y(
        n2471) );
  INV U3865 ( .A(n3490), .Y(n3489) );
  AOI222 U3866 ( .A0(n2655), .A1(\uut/mult_mant/c1 [7]), .B0(n2653), .B1(
        \uut/mult_mant/b1 [7]), .C0(n2661), .C1(\uut/mult_mant/a1 [7]), .Y(
        n3490) );
  OAI2BB1 U3867 ( .A0N(n3465), .A1N(n2540), .B0(n3491), .Y(n3476) );
  OAI2BB2 U3868 ( .B0(n3492), .B1(n3466), .A0N(n2541), .A1N(n3493), .Y(n3475)
         );
  INV U3869 ( .A(n3469), .Y(n3493) );
  INV U3870 ( .A(n3465), .Y(n3466) );
  INV U3871 ( .A(n3460), .Y(n3492) );
  NOR2B U3872 ( .AN(n2541), .B(n3452), .Y(n3460) );
  OAI2BB2 U3873 ( .B0(n2541), .B1(n3469), .A0N(n3465), .A1N(n3453), .Y(n3474)
         );
  NOR2B U3874 ( .AN(n2541), .B(\uut/mult_mant/mult8_cnt[1] ), .Y(n3453) );
  NAND2B U3875 ( .AN(\uut/mult_mant/mult8_cnt[2] ), .B(n3458), .Y(n3469) );
  INV U3876 ( .A(\uut/mult_mant/mult8_cnt[3] ), .Y(n3458) );
  MX2 U3877 ( .A(\uut/mult_mant/in2_segment [0]), .B(n3494), .S0(n2783), .Y(
        n2470) );
  INV U3878 ( .A(n3495), .Y(n3494) );
  AOI222 U3879 ( .A0(n2663), .A1(\uut/mult_mant/a2 [0]), .B0(
        \uut/mult_mant/b2 [0]), .B1(n2713), .C0(\uut/mult_mant/c2 [0]), .C1(
        n2718), .Y(n3495) );
  MX2 U3880 ( .A(\uut/mult_mant/in2_segment [1]), .B(n3497), .S0(n2783), .Y(
        n2469) );
  INV U3881 ( .A(n3498), .Y(n3497) );
  AOI222 U3882 ( .A0(n2663), .A1(\uut/mult_mant/a2 [1]), .B0(
        \uut/mult_mant/b2 [1]), .B1(n2713), .C0(\uut/mult_mant/c2 [1]), .C1(
        n2718), .Y(n3498) );
  MX2 U3883 ( .A(\uut/mult_mant/in2_segment [2]), .B(n3499), .S0(n2783), .Y(
        n2468) );
  INV U3884 ( .A(n3500), .Y(n3499) );
  AOI222 U3885 ( .A0(n2663), .A1(\uut/mult_mant/a2 [2]), .B0(
        \uut/mult_mant/b2 [2]), .B1(n2713), .C0(\uut/mult_mant/c2 [2]), .C1(
        n2718), .Y(n3500) );
  MX2 U3886 ( .A(\uut/mult_mant/in2_segment [3]), .B(n3501), .S0(n3471), .Y(
        n2467) );
  INV U3887 ( .A(n3502), .Y(n3501) );
  AOI222 U3888 ( .A0(n2663), .A1(\uut/mult_mant/a2 [3]), .B0(n2713), .B1(
        \uut/mult_mant/b2 [3]), .C0(\uut/mult_mant/c2 [3]), .C1(n2718), .Y(
        n3502) );
  MX2 U3889 ( .A(\uut/mult_mant/in2_segment [4]), .B(n3503), .S0(n2783), .Y(
        n2466) );
  INV U3890 ( .A(n3504), .Y(n3503) );
  AOI222 U3891 ( .A0(n2663), .A1(\uut/mult_mant/a2 [4]), .B0(n2713), .B1(
        \uut/mult_mant/b2 [4]), .C0(\uut/mult_mant/c2 [4]), .C1(n2718), .Y(
        n3504) );
  MX2 U3892 ( .A(\uut/mult_mant/in2_segment [5]), .B(n3505), .S0(n3471), .Y(
        n2465) );
  INV U3893 ( .A(n3506), .Y(n3505) );
  AOI222 U3894 ( .A0(n2663), .A1(\uut/mult_mant/a2 [5]), .B0(n2713), .B1(
        \uut/mult_mant/b2 [5]), .C0(\uut/mult_mant/c2 [5]), .C1(n2718), .Y(
        n3506) );
  MX2 U3895 ( .A(\uut/mult_mant/in2_segment [6]), .B(n3507), .S0(n2783), .Y(
        n2464) );
  INV U3896 ( .A(n3508), .Y(n3507) );
  AOI222 U3897 ( .A0(n2663), .A1(\uut/mult_mant/a2 [6]), .B0(n2713), .B1(
        \uut/mult_mant/b2 [6]), .C0(\uut/mult_mant/c2 [6]), .C1(n2718), .Y(
        n3508) );
  MX2 U3898 ( .A(\uut/mult_mant/in2_segment [7]), .B(n3509), .S0(n3471), .Y(
        n2463) );
  NOR2B U3899 ( .AN(n2697), .B(n2784), .Y(n3471) );
  OAI2BB2 U3900 ( .B0(n3510), .B1(n3511), .A0N(n3512), .A1N(
        \uut/mult_mant/mult8_cnt[3] ), .Y(n2784) );
  NOR2B U3901 ( .AN(rst_n), .B(n3513), .Y(n3511) );
  NOR2 U3902 ( .A(n2528), .B(\uut/mult_mant/mult_end [3]), .Y(n3513) );
  NOR2 U3903 ( .A(n3512), .B(\uut/mult_mant/mult8_cnt[3] ), .Y(n3510) );
  NOR2 U3904 ( .A(n3514), .B(n3515), .Y(n3512) );
  NOR2B U3905 ( .AN(n3516), .B(\uut/mult_mant/mult8_cnt[2] ), .Y(n3515) );
  NOR4BB U3906 ( .AN(rst_n), .BN(\uut/mult_mant/mult_end [2]), .C(n3517), .D(
        n2696), .Y(n3514) );
  NOR2B U3907 ( .AN(\uut/mult_mant/mult8_cnt[2] ), .B(n3516), .Y(n3517) );
  AOI211 U3908 ( .A0(n3518), .A1(n2697), .B0(\uut/mult_mant/mult8_cnt[1] ), 
        .C0(n2541), .Y(n3516) );
  NOR2B U3909 ( .AN(rst_n), .B(\uut/mult_mant/mult_end [3]), .Y(n3518) );
  NOR3B U3910 ( .AN(\uut/mult_mant/state[0] ), .B(\uut/mult_mant/state[2] ), 
        .C(\uut/mult_mant/state[1] ), .Y(n2785) );
  INV U3911 ( .A(n3519), .Y(n3509) );
  AOI222 U3912 ( .A0(n2663), .A1(\uut/mult_mant/a2 [7]), .B0(n2713), .B1(
        \uut/mult_mant/b2 [7]), .C0(\uut/mult_mant/c2 [7]), .C1(n2718), .Y(
        n3519) );
  INV U3913 ( .A(\uut/mult_mant/mult8_cnt[1] ), .Y(n3452) );
  NOR2B U3914 ( .AN(\uut/mult_mant/mult8_cnt[2] ), .B(n2540), .Y(n3520) );
  OAI2BB1 U3915 ( .A0N(n3465), .A1N(n2541), .B0(n3491), .Y(n3496) );
  INV U3916 ( .A(n3470), .Y(n3491) );
  NOR4B U3917 ( .AN(\uut/mult_mant/mult8_cnt[3] ), .B(
        \uut/mult_mant/mult8_cnt[1] ), .C(n2541), .D(
        \uut/mult_mant/mult8_cnt[2] ), .Y(n3470) );
  NOR2B U3918 ( .AN(\uut/mult_mant/mult8_cnt[2] ), .B(
        \uut/mult_mant/mult8_cnt[3] ), .Y(n3465) );
  OAI31 U3919 ( .A0(n2787), .A1(n2641), .A2(n2878), .B0(n3521), .Y(n2462) );
  INV U3920 ( .A(n3392), .Y(n3521) );
  NOR2B U3921 ( .AN(n3522), .B(n2640), .Y(n3392) );
  MX2 U3922 ( .A(\uut/mult_mant/temp_product[21] ), .B(
        \uut/mult_mant/temp_product[47] ), .S0(data_type), .Y(n3522) );
  INV U3923 ( .A(\uut/normalize ), .Y(n2878) );
  MX2 U3924 ( .A(n3523), .B(n3524), .S0(n2641), .Y(n2461) );
  NOR3B U3925 ( .AN(\uut/mult_mant/state[0] ), .B(\uut/mult_mant/state[2] ), 
        .C(n3525), .Y(n4988) );
  INV U3926 ( .A(\uut/mult_mant/state[1] ), .Y(n3525) );
  MX2 U3927 ( .A(\uut/mult_mant/temp_product[20] ), .B(
        \uut/mult_mant/temp_product[46] ), .S0(data_type), .Y(n3524) );
  NOR2B U3928 ( .AN(\uut/more_than_1 ), .B(n2787), .Y(n3523) );
  NOR2B U3929 ( .AN(n3391), .B(\uut/mult_mant/state[1] ), .Y(n2787) );
  NOR2 U3930 ( .A(\uut/mult_mant/state[0] ), .B(\uut/mult_mant/state[2] ), .Y(
        n3391) );
  OAI2BB1 U3931 ( .A0N(\uut/in1_32_reg[31] ), .A1N(n2738), .B0(n3526), .Y(
        n2400) );
  OAI2BB1 U3932 ( .A0N(\uut/in1_32_reg[30] ), .A1N(n2739), .B0(n3527), .Y(
        n2399) );
  OAI2BB1 U3933 ( .A0N(\uut/in1_32_reg[29] ), .A1N(n2738), .B0(n3528), .Y(
        n2398) );
  OAI2BB1 U3934 ( .A0N(\uut/in1_32_reg[28] ), .A1N(n2739), .B0(n3529), .Y(
        n2397) );
  OAI21 U3935 ( .A0(n2776), .A1(n3530), .B0(n3531), .Y(n2396) );
  OAI21 U3936 ( .A0(n2774), .A1(n3532), .B0(n3533), .Y(n2395) );
  OAI21 U3937 ( .A0(n2776), .A1(n3534), .B0(n3535), .Y(n2394) );
  OAI2BB1 U3938 ( .A0N(\uut/in1_32_reg[24] ), .A1N(n2738), .B0(n3536), .Y(
        n2393) );
  OAI21 U3939 ( .A0(n2776), .A1(n3537), .B0(n3538), .Y(n2392) );
  OAI21 U3940 ( .A0(n2529), .A1(n3539), .B0(n3540), .Y(n2391) );
  OAI21 U3941 ( .A0(n2776), .A1(n3541), .B0(n3542), .Y(n2390) );
  OAI21 U3942 ( .A0(n2775), .A1(n3543), .B0(n3544), .Y(n2389) );
  OAI21 U3943 ( .A0(n2775), .A1(n3545), .B0(n3546), .Y(n2388) );
  OAI21 U3944 ( .A0(n2529), .A1(n3547), .B0(n3548), .Y(n2387) );
  OAI21 U3945 ( .A0(n2775), .A1(n3549), .B0(n3550), .Y(n2386) );
  OAI21 U3946 ( .A0(n2773), .A1(n3551), .B0(n3552), .Y(n2385) );
  MX2 U3947 ( .A(\uut/in1_32_reg[15] ), .B(in1_disp[15]), .S0(n2529), .Y(n2384) );
  MX2 U3948 ( .A(\uut/in1_32_reg[14] ), .B(n2629), .S0(n2773), .Y(n2383) );
  MX2 U3949 ( .A(\uut/in1_32_reg[13] ), .B(in1_disp[13]), .S0(n2773), .Y(n2382) );
  MX2 U3950 ( .A(\uut/in1_32_reg[12] ), .B(n2627), .S0(n2773), .Y(n2381) );
  MX2 U3951 ( .A(\uut/in1_32_reg[11] ), .B(in1_disp[11]), .S0(n2773), .Y(n2380) );
  MX2 U3952 ( .A(\uut/in1_32_reg[10] ), .B(in1_disp[10]), .S0(n2774), .Y(n2379) );
  MX2 U3953 ( .A(\uut/in1_32_reg[9] ), .B(in1_disp[9]), .S0(n2774), .Y(n2378)
         );
  MX2 U3954 ( .A(\uut/in1_32_reg[8] ), .B(in1_disp[8]), .S0(n2774), .Y(n2377)
         );
  MX2 U3955 ( .A(\uut/in1_32_reg[7] ), .B(in1_disp[7]), .S0(n2529), .Y(n2376)
         );
  MX2 U3956 ( .A(\uut/in1_32_reg[6] ), .B(n2633), .S0(n2776), .Y(n2375) );
  MX2 U3957 ( .A(\uut/in1_32_reg[5] ), .B(in1_disp[5]), .S0(n2776), .Y(n2374)
         );
  MX2 U3958 ( .A(\uut/in1_32_reg[4] ), .B(n2631), .S0(n2776), .Y(n2373) );
  MX2 U3959 ( .A(\uut/in1_32_reg[3] ), .B(in1_disp[3]), .S0(n2529), .Y(n2372)
         );
  MX2 U3960 ( .A(\uut/in1_32_reg[2] ), .B(n2637), .S0(n2775), .Y(n2371) );
  MX2 U3961 ( .A(\uut/in1_32_reg[1] ), .B(in1_disp[1]), .S0(n2775), .Y(n2370)
         );
  MX2 U3962 ( .A(\uut/in1_32_reg[0] ), .B(n2635), .S0(n2775), .Y(n2369) );
  OAI2BB1 U3963 ( .A0N(\uut/in2_32_reg[31] ), .A1N(n2739), .B0(n3553), .Y(
        n2368) );
  OAI2BB1 U3964 ( .A0N(\uut/in2_32_reg[30] ), .A1N(n2738), .B0(n3554), .Y(
        n2367) );
  OAI2BB1 U3965 ( .A0N(\uut/in2_32_reg[29] ), .A1N(n2739), .B0(n3555), .Y(
        n2366) );
  OAI2BB1 U3966 ( .A0N(\uut/in2_32_reg[28] ), .A1N(n2738), .B0(n3556), .Y(
        n2365) );
  OAI21 U3967 ( .A0(n2773), .A1(n3557), .B0(n3558), .Y(n2364) );
  OAI21 U3968 ( .A0(n2529), .A1(n3559), .B0(n3560), .Y(n2363) );
  OAI21 U3969 ( .A0(n2773), .A1(n3561), .B0(n3562), .Y(n2362) );
  OAI2BB1 U3970 ( .A0N(\uut/in2_32_reg[24] ), .A1N(n2739), .B0(n3563), .Y(
        n2361) );
  OAI21 U3971 ( .A0(n2774), .A1(n3564), .B0(n3565), .Y(n2360) );
  OAI21 U3972 ( .A0(n2774), .A1(n3566), .B0(n3567), .Y(n2359) );
  OAI21 U3973 ( .A0(n2774), .A1(n3568), .B0(n3569), .Y(n2358) );
  OAI21 U3974 ( .A0(n2774), .A1(n3570), .B0(n3571), .Y(n2357) );
  OAI21 U3975 ( .A0(n2776), .A1(n3572), .B0(n3573), .Y(n2356) );
  OAI21 U3976 ( .A0(n2776), .A1(n3574), .B0(n3575), .Y(n2355) );
  OAI21 U3977 ( .A0(n2529), .A1(n3576), .B0(n3577), .Y(n2354) );
  OAI21 U3978 ( .A0(n2776), .A1(n3578), .B0(n3579), .Y(n2353) );
  MX2 U3979 ( .A(\uut/in2_32_reg[15] ), .B(in2_disp[15]), .S0(n2529), .Y(n2352) );
  MX2 U3980 ( .A(\uut/in2_32_reg[14] ), .B(n2609), .S0(n2773), .Y(n2351) );
  MX2 U3981 ( .A(\uut/in2_32_reg[13] ), .B(in2_disp[13]), .S0(n2773), .Y(n2350) );
  MX2 U3982 ( .A(\uut/in2_32_reg[12] ), .B(n2607), .S0(n2773), .Y(n2349) );
  MX2 U3983 ( .A(\uut/in2_32_reg[11] ), .B(in2_disp[11]), .S0(n2529), .Y(n2348) );
  MX2 U3984 ( .A(\uut/in2_32_reg[10] ), .B(in2_disp[10]), .S0(n2774), .Y(n2347) );
  MX2 U3985 ( .A(\uut/in2_32_reg[9] ), .B(in2_disp[9]), .S0(n2774), .Y(n2346)
         );
  MX2 U3986 ( .A(\uut/in2_32_reg[8] ), .B(in2_disp[8]), .S0(n2774), .Y(n2345)
         );
  MX2 U3987 ( .A(\uut/in2_32_reg[7] ), .B(in2_disp[7]), .S0(n2529), .Y(n2344)
         );
  MX2 U3988 ( .A(\uut/in2_32_reg[6] ), .B(n2613), .S0(n2776), .Y(n2343) );
  MX2 U3989 ( .A(\uut/in2_32_reg[5] ), .B(in2_disp[5]), .S0(n2776), .Y(n2342)
         );
  MX2 U3990 ( .A(\uut/in2_32_reg[4] ), .B(n2611), .S0(n2776), .Y(n2341) );
  MX2 U3991 ( .A(\uut/in2_32_reg[3] ), .B(in2_disp[3]), .S0(n2529), .Y(n2340)
         );
  MX2 U3992 ( .A(\uut/in2_32_reg[2] ), .B(n2617), .S0(n2775), .Y(n2339) );
  MX2 U3993 ( .A(\uut/in2_32_reg[1] ), .B(in2_disp[1]), .S0(n2775), .Y(n2338)
         );
  MX2 U3994 ( .A(\uut/in2_32_reg[0] ), .B(n2615), .S0(n2775), .Y(n2337) );
  OAI2BB1 U3995 ( .A0N(\uut/in1_16_reg[15] ), .A1N(n2738), .B0(n3526), .Y(
        n2336) );
  NAND2 U3996 ( .A(n2775), .B(n2619), .Y(n3526) );
  OAI2BB1 U3997 ( .A0N(\uut/in1_16_reg[14] ), .A1N(n2739), .B0(n3527), .Y(
        n2335) );
  NAND2 U3998 ( .A(n2775), .B(in1_disp[30]), .Y(n3527) );
  OAI21 U3999 ( .A0(n2773), .A1(n3580), .B0(n3528), .Y(n2334) );
  NAND2 U4000 ( .A(n2775), .B(in1_disp[29]), .Y(n3528) );
  OAI21 U4001 ( .A0(n2773), .A1(n3581), .B0(n3529), .Y(n2333) );
  NAND2 U4002 ( .A(n2773), .B(n2679), .Y(n3529) );
  OAI2BB1 U4003 ( .A0N(\uut/in1_16_reg[11] ), .A1N(n2738), .B0(n3531), .Y(
        n2332) );
  NAND2 U4004 ( .A(n2529), .B(n2621), .Y(n3531) );
  OAI21 U4005 ( .A0(n2773), .A1(n3582), .B0(n3533), .Y(n2331) );
  NAND2 U4006 ( .A(n2776), .B(in1_disp[26]), .Y(n3533) );
  OAI2BB1 U4007 ( .A0N(\uut/in1_16_reg[9] ), .A1N(n2739), .B0(n3535), .Y(n2330) );
  NAND2 U4008 ( .A(n2774), .B(in1_disp[25]), .Y(n3535) );
  OAI2BB1 U4009 ( .A0N(\uut/in1_16_reg[8] ), .A1N(n2738), .B0(n3536), .Y(n2329) );
  NAND2 U4010 ( .A(n2776), .B(in1_disp[24]), .Y(n3536) );
  OAI2BB1 U4011 ( .A0N(\uut/in1_16_reg[7] ), .A1N(n2739), .B0(n3538), .Y(n2328) );
  NAND2 U4012 ( .A(n2774), .B(n2623), .Y(n3538) );
  OAI2BB1 U4013 ( .A0N(\uut/in1_16_reg[6] ), .A1N(n2738), .B0(n3540), .Y(n2327) );
  NAND2 U4014 ( .A(n2774), .B(in1_disp[22]), .Y(n3540) );
  OAI2BB1 U4015 ( .A0N(\uut/in1_16_reg[5] ), .A1N(n2739), .B0(n3542), .Y(n2326) );
  NAND2 U4016 ( .A(n2774), .B(in1_disp[21]), .Y(n3542) );
  OAI2BB1 U4017 ( .A0N(\uut/in1_16_reg[4] ), .A1N(n2738), .B0(n3544), .Y(n2325) );
  NAND2 U4018 ( .A(n2529), .B(n2673), .Y(n3544) );
  OAI2BB1 U4019 ( .A0N(\uut/in1_16_reg[3] ), .A1N(n2739), .B0(n3546), .Y(n2324) );
  NAND2 U4020 ( .A(n2776), .B(n2625), .Y(n3546) );
  OAI2BB1 U4021 ( .A0N(\uut/in1_16_reg[2] ), .A1N(n2738), .B0(n3548), .Y(n2323) );
  NAND2 U4022 ( .A(n2776), .B(in1_disp[18]), .Y(n3548) );
  OAI2BB1 U4023 ( .A0N(\uut/in1_16_reg[1] ), .A1N(n2739), .B0(n3550), .Y(n2322) );
  NAND2 U4024 ( .A(n2776), .B(in1_disp[17]), .Y(n3550) );
  OAI2BB1 U4025 ( .A0N(\uut/in1_16_reg[0] ), .A1N(n2738), .B0(n3552), .Y(n2321) );
  NAND2 U4026 ( .A(n2774), .B(n2675), .Y(n3552) );
  OAI2BB1 U4027 ( .A0N(\uut/in2_16_reg[15] ), .A1N(n2739), .B0(n3553), .Y(
        n2320) );
  NAND2 U4028 ( .A(n2775), .B(n2599), .Y(n3553) );
  OAI2BB1 U4029 ( .A0N(\uut/in2_16_reg[14] ), .A1N(n2738), .B0(n3554), .Y(
        n2319) );
  NAND2 U4030 ( .A(n2775), .B(in2_disp[30]), .Y(n3554) );
  OAI21 U4031 ( .A0(n2776), .A1(n3583), .B0(n3555), .Y(n2318) );
  NAND2 U4032 ( .A(n2529), .B(in2_disp[29]), .Y(n3555) );
  OAI21 U4033 ( .A0(n2773), .A1(n3584), .B0(n3556), .Y(n2317) );
  NAND2 U4034 ( .A(n2775), .B(n2681), .Y(n3556) );
  OAI2BB1 U4035 ( .A0N(\uut/in2_16_reg[11] ), .A1N(n2739), .B0(n3558), .Y(
        n2316) );
  NAND2 U4036 ( .A(n2775), .B(n2601), .Y(n3558) );
  OAI21 U4037 ( .A0(n2775), .A1(n3585), .B0(n3560), .Y(n2315) );
  NAND2 U4038 ( .A(n2774), .B(in2_disp[26]), .Y(n3560) );
  OAI2BB1 U4039 ( .A0N(\uut/in2_16_reg[9] ), .A1N(n2738), .B0(n3562), .Y(n2314) );
  NAND2 U4040 ( .A(n2775), .B(in2_disp[25]), .Y(n3562) );
  OAI2BB1 U4041 ( .A0N(\uut/in2_16_reg[8] ), .A1N(n2739), .B0(n3563), .Y(n2313) );
  NAND2 U4042 ( .A(n2773), .B(in2_disp[24]), .Y(n3563) );
  OAI2BB1 U4043 ( .A0N(\uut/in2_16_reg[7] ), .A1N(n2738), .B0(n3565), .Y(n2312) );
  NAND2 U4044 ( .A(n2529), .B(n2603), .Y(n3565) );
  OAI2BB1 U4045 ( .A0N(\uut/in2_16_reg[6] ), .A1N(n2739), .B0(n3567), .Y(n2311) );
  NAND2 U4046 ( .A(n2776), .B(in2_disp[22]), .Y(n3567) );
  OAI2BB1 U4047 ( .A0N(\uut/in2_16_reg[5] ), .A1N(n2738), .B0(n3569), .Y(n2310) );
  NAND2 U4048 ( .A(n2773), .B(in2_disp[21]), .Y(n3569) );
  OAI2BB1 U4049 ( .A0N(\uut/in2_16_reg[4] ), .A1N(n2739), .B0(n3571), .Y(n2309) );
  NAND2 U4050 ( .A(n2773), .B(n2683), .Y(n3571) );
  OAI2BB1 U4051 ( .A0N(\uut/in2_16_reg[3] ), .A1N(n2738), .B0(n3573), .Y(n2308) );
  NAND2 U4052 ( .A(n2773), .B(n2605), .Y(n3573) );
  OAI2BB1 U4053 ( .A0N(\uut/in2_16_reg[2] ), .A1N(n2739), .B0(n3575), .Y(n2307) );
  NAND2 U4054 ( .A(n2775), .B(in2_disp[18]), .Y(n3575) );
  OAI2BB1 U4055 ( .A0N(\uut/in2_16_reg[1] ), .A1N(n2738), .B0(n3577), .Y(n2306) );
  NAND2 U4056 ( .A(n2774), .B(in2_disp[17]), .Y(n3577) );
  OAI2BB1 U4057 ( .A0N(\uut/in2_16_reg[0] ), .A1N(n2739), .B0(n3579), .Y(n2305) );
  NAND2 U4058 ( .A(n2774), .B(n2677), .Y(n3579) );
  OAI2BB2 U4059 ( .B0(n2545), .B1(n3586), .A0N(\uut/mult_mant/b1 [3]), .A1N(
        n2766), .Y(n2293) );
  INV U4060 ( .A(\uut/in1_32_reg[11] ), .Y(n3586) );
  OAI2BB2 U4061 ( .B0(n2544), .B1(n3587), .A0N(\uut/mult_mant/b1 [4]), .A1N(
        n2768), .Y(n2292) );
  INV U4062 ( .A(\uut/in1_32_reg[12] ), .Y(n3587) );
  OAI2BB2 U4063 ( .B0(n2545), .B1(n3588), .A0N(\uut/mult_mant/b1 [5]), .A1N(
        n2767), .Y(n2291) );
  INV U4064 ( .A(\uut/in1_32_reg[13] ), .Y(n3588) );
  OAI2BB2 U4065 ( .B0(n2544), .B1(n3589), .A0N(\uut/mult_mant/b1 [6]), .A1N(
        n2766), .Y(n2290) );
  INV U4066 ( .A(\uut/in1_32_reg[14] ), .Y(n3589) );
  OAI2BB2 U4067 ( .B0(n2545), .B1(n3590), .A0N(\uut/mult_mant/b1 [7]), .A1N(
        n2768), .Y(n2289) );
  INV U4068 ( .A(\uut/in1_32_reg[15] ), .Y(n3590) );
  OAI2BB2 U4069 ( .B0(n2544), .B1(n3551), .A0N(\uut/mult_mant/a1 [0]), .A1N(
        n2767), .Y(n2288) );
  INV U4070 ( .A(\uut/in1_32_reg[16] ), .Y(n3551) );
  OAI2BB2 U4071 ( .B0(n2545), .B1(n3549), .A0N(\uut/mult_mant/a1 [1]), .A1N(
        n2766), .Y(n2287) );
  INV U4072 ( .A(\uut/in1_32_reg[17] ), .Y(n3549) );
  OAI2BB2 U4073 ( .B0(n2544), .B1(n3547), .A0N(\uut/mult_mant/a1 [2]), .A1N(
        n2768), .Y(n2286) );
  INV U4074 ( .A(\uut/in1_32_reg[18] ), .Y(n3547) );
  OAI2BB2 U4075 ( .B0(n2545), .B1(n3545), .A0N(\uut/mult_mant/a1 [3]), .A1N(
        n2767), .Y(n2285) );
  INV U4076 ( .A(\uut/in1_32_reg[19] ), .Y(n3545) );
  OAI2BB2 U4077 ( .B0(n2544), .B1(n3543), .A0N(\uut/mult_mant/a1 [4]), .A1N(
        n2766), .Y(n2284) );
  INV U4078 ( .A(\uut/in1_32_reg[20] ), .Y(n3543) );
  OAI2BB2 U4079 ( .B0(n2545), .B1(n3541), .A0N(\uut/mult_mant/a1 [5]), .A1N(
        n2768), .Y(n2283) );
  INV U4080 ( .A(\uut/in1_32_reg[21] ), .Y(n3541) );
  OAI2BB2 U4081 ( .B0(n2544), .B1(n3539), .A0N(\uut/mult_mant/a1 [6]), .A1N(
        n2767), .Y(n2282) );
  INV U4082 ( .A(\uut/in1_32_reg[22] ), .Y(n3539) );
  OAI2BB2 U4083 ( .B0(n2533), .B1(n2545), .A0N(\uut/mult_mant/a1 [7]), .A1N(
        n2766), .Y(n2281) );
  NOR4BB U4084 ( .AN(n3591), .BN(n3592), .C(n2922), .D(n3593), .Y(n2858) );
  MX2 U4085 ( .A(n2537), .B(n3595), .S0(data_type), .Y(n3593) );
  MX2 U4086 ( .A(\uut/in1_16_reg[14] ), .B(\uut/in1_32_reg[27] ), .S0(
        data_type), .Y(n2922) );
  NOR2 U4087 ( .A(n2911), .B(n2907), .Y(n3592) );
  MX2 U4088 ( .A(\uut/in1_16_reg[13] ), .B(\uut/in1_32_reg[26] ), .S0(
        data_type), .Y(n2907) );
  MX2 U4089 ( .A(\uut/in1_16_reg[12] ), .B(\uut/in1_32_reg[25] ), .S0(
        data_type), .Y(n2911) );
  NOR4BB U4090 ( .AN(n3596), .BN(n2803), .C(n2898), .D(n2917), .Y(n3591) );
  NOR2B U4091 ( .AN(\uut/in1_32_reg[29] ), .B(n4961), .Y(n2917) );
  NOR2B U4092 ( .AN(\uut/in1_32_reg[28] ), .B(n4961), .Y(n2898) );
  NOR2 U4093 ( .A(n2912), .B(n2915), .Y(n3596) );
  MX2 U4094 ( .A(\uut/in1_16_reg[11] ), .B(\uut/in1_32_reg[24] ), .S0(
        data_type), .Y(n2915) );
  INV U4095 ( .A(n2924), .Y(n2912) );
  MX2 U4096 ( .A(n3582), .B(n3537), .S0(data_type), .Y(n2924) );
  OAI2BB2 U4097 ( .B0(n2544), .B1(n3597), .A0N(\uut/mult_mant/b2 [3]), .A1N(
        n2768), .Y(n2269) );
  INV U4098 ( .A(\uut/in2_32_reg[11] ), .Y(n3597) );
  OAI2BB2 U4099 ( .B0(n2545), .B1(n3598), .A0N(\uut/mult_mant/b2 [4]), .A1N(
        n2767), .Y(n2268) );
  INV U4100 ( .A(\uut/in2_32_reg[12] ), .Y(n3598) );
  OAI2BB2 U4101 ( .B0(n2544), .B1(n3599), .A0N(\uut/mult_mant/b2 [5]), .A1N(
        n2766), .Y(n2267) );
  INV U4102 ( .A(\uut/in2_32_reg[13] ), .Y(n3599) );
  OAI2BB2 U4103 ( .B0(n2545), .B1(n3600), .A0N(\uut/mult_mant/b2 [6]), .A1N(
        n2768), .Y(n2266) );
  INV U4104 ( .A(\uut/in2_32_reg[14] ), .Y(n3600) );
  OAI2BB2 U4105 ( .B0(n2544), .B1(n3601), .A0N(\uut/mult_mant/b2 [7]), .A1N(
        n2767), .Y(n2265) );
  INV U4106 ( .A(\uut/in2_32_reg[15] ), .Y(n3601) );
  OAI2BB2 U4107 ( .B0(n2545), .B1(n3578), .A0N(\uut/mult_mant/a2 [0]), .A1N(
        n2766), .Y(n2264) );
  INV U4108 ( .A(\uut/in2_32_reg[16] ), .Y(n3578) );
  OAI2BB2 U4109 ( .B0(n2544), .B1(n3576), .A0N(\uut/mult_mant/a2 [1]), .A1N(
        n2768), .Y(n2263) );
  INV U4110 ( .A(\uut/in2_32_reg[17] ), .Y(n3576) );
  OAI2BB2 U4111 ( .B0(n2545), .B1(n3574), .A0N(\uut/mult_mant/a2 [2]), .A1N(
        n2767), .Y(n2262) );
  INV U4112 ( .A(\uut/in2_32_reg[18] ), .Y(n3574) );
  OAI2BB2 U4113 ( .B0(n2544), .B1(n3572), .A0N(\uut/mult_mant/a2 [3]), .A1N(
        n2766), .Y(n2261) );
  INV U4114 ( .A(\uut/in2_32_reg[19] ), .Y(n3572) );
  OAI2BB2 U4115 ( .B0(n2545), .B1(n3570), .A0N(\uut/mult_mant/a2 [4]), .A1N(
        n2768), .Y(n2260) );
  INV U4116 ( .A(\uut/in2_32_reg[20] ), .Y(n3570) );
  OAI2BB2 U4117 ( .B0(n2544), .B1(n3568), .A0N(\uut/mult_mant/a2 [5]), .A1N(
        n2767), .Y(n2259) );
  INV U4118 ( .A(\uut/in2_32_reg[21] ), .Y(n3568) );
  OAI2BB2 U4119 ( .B0(n2545), .B1(n3566), .A0N(\uut/mult_mant/a2 [6]), .A1N(
        n2766), .Y(n2258) );
  INV U4120 ( .A(\uut/in2_32_reg[22] ), .Y(n3566) );
  OAI2BB2 U4121 ( .B0(n2870), .B1(n2544), .A0N(\uut/mult_mant/a2 [7]), .A1N(
        n2768), .Y(n2257) );
  INV U4122 ( .A(n2902), .Y(n2870) );
  AOI22 U4123 ( .A0(n3602), .A1(n3603), .B0(n3604), .B1(n2534), .Y(n2902) );
  OAI222 U4124 ( .A0(n3605), .A1(n3016), .B0(n3606), .B1(n2763), .C0(n3068), 
        .C1(n3608), .Y(n2256) );
  INV U4125 ( .A(\uut/mult_mant/temp_product[10] ), .Y(n3068) );
  INV U4126 ( .A(\uut/mant_out[0] ), .Y(n3606) );
  INV U4127 ( .A(\uut/mult_mant/temp_product[23] ), .Y(n3016) );
  OAI222 U4128 ( .A0(n3605), .A1(n3012), .B0(n3609), .B1(n2763), .C0(n3064), 
        .C1(n3608), .Y(n2255) );
  INV U4129 ( .A(\uut/mult_mant/temp_product[11] ), .Y(n3064) );
  INV U4130 ( .A(\uut/mult_mant/temp_product[24] ), .Y(n3012) );
  OAI222 U4131 ( .A0(n3605), .A1(n3008), .B0(n3610), .B1(n2763), .C0(n3060), 
        .C1(n3608), .Y(n2254) );
  INV U4132 ( .A(\uut/mult_mant/temp_product[12] ), .Y(n3060) );
  INV U4133 ( .A(\uut/mant_out[2] ), .Y(n3610) );
  INV U4134 ( .A(\uut/mult_mant/temp_product[25] ), .Y(n3008) );
  OAI222 U4135 ( .A0(n3605), .A1(n3004), .B0(n3611), .B1(n2763), .C0(n3056), 
        .C1(n3608), .Y(n2253) );
  INV U4136 ( .A(\uut/mult_mant/temp_product[13] ), .Y(n3056) );
  INV U4137 ( .A(\uut/mant_out[3] ), .Y(n3611) );
  INV U4138 ( .A(\uut/mult_mant/temp_product[26] ), .Y(n3004) );
  OAI222 U4139 ( .A0(n3605), .A1(n3000), .B0(n3612), .B1(n2763), .C0(n3052), 
        .C1(n3608), .Y(n2252) );
  INV U4140 ( .A(\uut/mult_mant/temp_product[14] ), .Y(n3052) );
  INV U4141 ( .A(\uut/mant_out[4] ), .Y(n3612) );
  INV U4142 ( .A(\uut/mult_mant/temp_product[27] ), .Y(n3000) );
  OAI222 U4143 ( .A0(n3605), .A1(n2996), .B0(n3613), .B1(n2763), .C0(n3048), 
        .C1(n3608), .Y(n2251) );
  INV U4144 ( .A(\uut/mult_mant/temp_product[15] ), .Y(n3048) );
  INV U4145 ( .A(\uut/mult_mant/temp_product[28] ), .Y(n2996) );
  OAI222 U4146 ( .A0(n3605), .A1(n2992), .B0(n3614), .B1(n2763), .C0(n3044), 
        .C1(n3608), .Y(n2250) );
  INV U4147 ( .A(\uut/mult_mant/temp_product[16] ), .Y(n3044) );
  INV U4148 ( .A(\uut/mant_out[6] ), .Y(n3614) );
  INV U4149 ( .A(\uut/mult_mant/temp_product[29] ), .Y(n2992) );
  OAI222 U4150 ( .A0(n3605), .A1(n2988), .B0(n3615), .B1(n2763), .C0(n3040), 
        .C1(n3608), .Y(n2249) );
  INV U4151 ( .A(\uut/mult_mant/temp_product[17] ), .Y(n3040) );
  INV U4152 ( .A(\uut/mant_out[7] ), .Y(n3615) );
  INV U4153 ( .A(\uut/mult_mant/temp_product[30] ), .Y(n2988) );
  OAI222 U4154 ( .A0(n3605), .A1(n2984), .B0(n3616), .B1(n2763), .C0(n3036), 
        .C1(n3608), .Y(n2248) );
  INV U4155 ( .A(\uut/mult_mant/temp_product[18] ), .Y(n3036) );
  INV U4156 ( .A(\uut/mant_out[8] ), .Y(n3616) );
  INV U4157 ( .A(\uut/mult_mant/temp_product[31] ), .Y(n2984) );
  OAI222 U4158 ( .A0(n3605), .A1(n2980), .B0(n3617), .B1(n2763), .C0(n3032), 
        .C1(n3608), .Y(n2247) );
  NAND2B U4159 ( .AN(data_type), .B(n2763), .Y(n3608) );
  INV U4160 ( .A(\uut/mult_mant/temp_product[19] ), .Y(n3032) );
  INV U4161 ( .A(\uut/mant_out[9] ), .Y(n3617) );
  INV U4162 ( .A(\uut/mult_mant/temp_product[32] ), .Y(n2980) );
  OAI2BB2 U4163 ( .B0(n2976), .B1(n3605), .A0N(\uut/mant_out[10] ), .A1N(n2762), .Y(n2246) );
  INV U4164 ( .A(\uut/mult_mant/temp_product[33] ), .Y(n2976) );
  OAI2BB2 U4165 ( .B0(n2972), .B1(n3605), .A0N(\uut/mant_out[11] ), .A1N(n2762), .Y(n2245) );
  INV U4166 ( .A(\uut/mult_mant/temp_product[34] ), .Y(n2972) );
  OAI2BB2 U4167 ( .B0(n2968), .B1(n3605), .A0N(\uut/mant_out[12] ), .A1N(n2762), .Y(n2244) );
  INV U4168 ( .A(\uut/mult_mant/temp_product[35] ), .Y(n2968) );
  OAI2BB2 U4169 ( .B0(n2964), .B1(n3605), .A0N(\uut/mant_out[13] ), .A1N(n2762), .Y(n2243) );
  INV U4170 ( .A(\uut/mult_mant/temp_product[36] ), .Y(n2964) );
  OAI2BB2 U4171 ( .B0(n2960), .B1(n3605), .A0N(\uut/mant_out[14] ), .A1N(n2762), .Y(n2242) );
  INV U4172 ( .A(\uut/mult_mant/temp_product[37] ), .Y(n2960) );
  OAI2BB2 U4173 ( .B0(n2956), .B1(n3605), .A0N(\uut/mant_out[15] ), .A1N(n2762), .Y(n2241) );
  INV U4174 ( .A(\uut/mult_mant/temp_product[38] ), .Y(n2956) );
  OAI2BB2 U4175 ( .B0(n2952), .B1(n3605), .A0N(\uut/mant_out[16] ), .A1N(n2762), .Y(n2240) );
  INV U4176 ( .A(\uut/mult_mant/temp_product[39] ), .Y(n2952) );
  OAI2BB2 U4177 ( .B0(n2948), .B1(n3605), .A0N(\uut/mant_out[17] ), .A1N(n2762), .Y(n2239) );
  INV U4178 ( .A(\uut/mult_mant/temp_product[40] ), .Y(n2948) );
  OAI2BB2 U4179 ( .B0(n2944), .B1(n3605), .A0N(\uut/mant_out[18] ), .A1N(n2762), .Y(n2238) );
  INV U4180 ( .A(\uut/mult_mant/temp_product[41] ), .Y(n2944) );
  OAI2BB2 U4181 ( .B0(n2940), .B1(n3605), .A0N(\uut/mant_out[19] ), .A1N(n2762), .Y(n2237) );
  INV U4182 ( .A(\uut/mult_mant/temp_product[42] ), .Y(n2940) );
  OAI2BB2 U4183 ( .B0(n2936), .B1(n3605), .A0N(\uut/mant_out[20] ), .A1N(n2762), .Y(n2236) );
  INV U4184 ( .A(\uut/mult_mant/temp_product[43] ), .Y(n2936) );
  OAI2BB2 U4185 ( .B0(n2932), .B1(n3605), .A0N(\uut/mant_out[21] ), .A1N(n2762), .Y(n2235) );
  INV U4186 ( .A(\uut/mult_mant/temp_product[44] ), .Y(n2932) );
  OAI2BB2 U4187 ( .B0(n2928), .B1(n3605), .A0N(\uut/mant_out[22] ), .A1N(n2762), .Y(n2234) );
  NAND2 U4188 ( .A(data_type), .B(n2763), .Y(n3605) );
  NOR3B U4189 ( .AN(\uut/mult_mant/state[2] ), .B(\uut/mult_mant/state[0] ), 
        .C(\uut/mult_mant/state[1] ), .Y(n3607) );
  INV U4190 ( .A(\uut/mult_mant/temp_product[45] ), .Y(n2928) );
  NAND4 U4191 ( .A(n3618), .B(n3619), .C(n3620), .D(n3621), .Y(disp2_seg[6])
         );
  AOI22 U4192 ( .A0(disp2_sel[6]), .A1(disp2_bit6[6]), .B0(disp2_sel[5]), .B1(
        disp2_bit5[6]), .Y(n3621) );
  AOI22 U4193 ( .A0(disp2_sel[4]), .A1(disp2_bit4[6]), .B0(disp2_sel[3]), .B1(
        disp2_bit3[6]), .Y(n3620) );
  AOI22 U4194 ( .A0(disp2_sel[2]), .A1(disp2_bit2[6]), .B0(disp2_sel[1]), .B1(
        disp2_bit1[6]), .Y(n3619) );
  AOI22 U4195 ( .A0(disp2_sel[7]), .A1(disp2_bit7[6]), .B0(disp2_sel[0]), .B1(
        disp2_bit0[6]), .Y(n3618) );
  NAND4 U4196 ( .A(n3622), .B(n3623), .C(n3624), .D(n3625), .Y(disp2_seg[5])
         );
  AOI22 U4197 ( .A0(disp2_sel[6]), .A1(disp2_bit6[5]), .B0(disp2_sel[5]), .B1(
        disp2_bit5[5]), .Y(n3625) );
  AOI22 U4198 ( .A0(disp2_sel[4]), .A1(disp2_bit4[5]), .B0(disp2_sel[3]), .B1(
        disp2_bit3[5]), .Y(n3624) );
  AOI22 U4199 ( .A0(disp2_sel[2]), .A1(disp2_bit2[5]), .B0(disp2_sel[1]), .B1(
        disp2_bit1[5]), .Y(n3623) );
  AOI22 U4200 ( .A0(disp2_sel[7]), .A1(disp2_bit7[5]), .B0(disp2_sel[0]), .B1(
        disp2_bit0[5]), .Y(n3622) );
  NAND4 U4201 ( .A(n3626), .B(n3627), .C(n3628), .D(n3629), .Y(disp2_seg[4])
         );
  AOI22 U4202 ( .A0(disp2_sel[6]), .A1(disp2_bit6[4]), .B0(disp2_sel[5]), .B1(
        disp2_bit5[4]), .Y(n3629) );
  AOI22 U4203 ( .A0(disp2_sel[4]), .A1(disp2_bit4[4]), .B0(disp2_sel[3]), .B1(
        disp2_bit3[4]), .Y(n3628) );
  AOI22 U4204 ( .A0(disp2_sel[2]), .A1(disp2_bit2[4]), .B0(disp2_sel[1]), .B1(
        disp2_bit1[4]), .Y(n3627) );
  AOI22 U4205 ( .A0(disp2_sel[7]), .A1(disp2_bit7[4]), .B0(disp2_sel[0]), .B1(
        disp2_bit0[4]), .Y(n3626) );
  NAND4 U4206 ( .A(n3630), .B(n3631), .C(n3632), .D(n3633), .Y(disp2_seg[3])
         );
  AOI22 U4207 ( .A0(disp2_sel[6]), .A1(disp2_bit6[3]), .B0(disp2_sel[5]), .B1(
        disp2_bit5[3]), .Y(n3633) );
  AOI22 U4208 ( .A0(disp2_sel[4]), .A1(disp2_bit4[3]), .B0(disp2_sel[3]), .B1(
        disp2_bit3[3]), .Y(n3632) );
  AOI22 U4209 ( .A0(disp2_sel[2]), .A1(disp2_bit2[3]), .B0(disp2_sel[1]), .B1(
        disp2_bit1[3]), .Y(n3631) );
  AOI22 U4210 ( .A0(disp2_sel[7]), .A1(disp2_bit7[3]), .B0(disp2_sel[0]), .B1(
        disp2_bit0[3]), .Y(n3630) );
  NAND4 U4211 ( .A(n3634), .B(n3635), .C(n3636), .D(n3637), .Y(disp2_seg[2])
         );
  AOI22 U4212 ( .A0(disp2_sel[6]), .A1(disp2_bit6[2]), .B0(disp2_sel[5]), .B1(
        disp2_bit5[2]), .Y(n3637) );
  AOI22 U4213 ( .A0(disp2_sel[4]), .A1(disp2_bit4[2]), .B0(disp2_sel[3]), .B1(
        disp2_bit3[2]), .Y(n3636) );
  AOI22 U4214 ( .A0(disp2_sel[2]), .A1(disp2_bit2[2]), .B0(disp2_sel[1]), .B1(
        disp2_bit1[2]), .Y(n3635) );
  AOI22 U4215 ( .A0(disp2_sel[7]), .A1(disp2_bit7[2]), .B0(disp2_sel[0]), .B1(
        disp2_bit0[2]), .Y(n3634) );
  NAND4 U4216 ( .A(n3638), .B(n3639), .C(n3640), .D(n3641), .Y(disp2_seg[1])
         );
  AOI22 U4217 ( .A0(disp2_sel[6]), .A1(disp2_bit6[1]), .B0(disp2_sel[5]), .B1(
        disp2_bit5[1]), .Y(n3641) );
  AOI22 U4218 ( .A0(disp2_sel[4]), .A1(disp2_bit4[1]), .B0(disp2_sel[3]), .B1(
        disp2_bit3[1]), .Y(n3640) );
  AOI22 U4219 ( .A0(disp2_sel[2]), .A1(disp2_bit2[1]), .B0(disp2_sel[1]), .B1(
        disp2_bit1[1]), .Y(n3639) );
  AOI22 U4220 ( .A0(disp2_sel[7]), .A1(disp2_bit7[1]), .B0(disp2_sel[0]), .B1(
        disp2_bit0[1]), .Y(n3638) );
  NAND4 U4221 ( .A(n3642), .B(n3643), .C(n3644), .D(n3645), .Y(disp2_seg[0])
         );
  AOI22 U4222 ( .A0(disp2_sel[6]), .A1(disp2_bit6[0]), .B0(disp2_sel[5]), .B1(
        disp2_bit5[0]), .Y(n3645) );
  NOR2B U4223 ( .AN(n3646), .B(n4979), .Y(n4996) );
  NOR2B U4224 ( .AN(n3647), .B(n3648), .Y(n4995) );
  AOI22 U4225 ( .A0(disp2_sel[4]), .A1(disp2_bit4[0]), .B0(disp2_sel[3]), .B1(
        disp2_bit3[0]), .Y(n3644) );
  NOR2B U4226 ( .AN(n3646), .B(disp2_sel_cnt[0]), .Y(n4997) );
  AOI22 U4227 ( .A0(disp2_sel[2]), .A1(disp2_bit2[0]), .B0(disp2_sel[1]), .B1(
        disp2_bit1[0]), .Y(n3643) );
  NOR2B U4228 ( .AN(n3649), .B(n4979), .Y(n5000) );
  NOR2B U4229 ( .AN(n3647), .B(disp2_sel_cnt[2]), .Y(n4999) );
  AOI22 U4230 ( .A0(disp2_sel[7]), .A1(disp2_bit7[0]), .B0(disp2_sel[0]), .B1(
        disp2_bit0[0]), .Y(n3642) );
  NAND4 U4231 ( .A(n3650), .B(n3651), .C(n3652), .D(n3653), .Y(disp1_seg[6])
         );
  AOI22 U4232 ( .A0(disp1_sel[6]), .A1(disp1_bit6[6]), .B0(disp1_sel[5]), .B1(
        disp1_bit5[6]), .Y(n3653) );
  AOI22 U4233 ( .A0(disp1_sel[4]), .A1(disp1_bit4[6]), .B0(disp1_sel[3]), .B1(
        disp1_bit3[6]), .Y(n3652) );
  AOI22 U4234 ( .A0(disp1_sel[2]), .A1(disp1_bit2[6]), .B0(disp1_sel[1]), .B1(
        disp1_bit1[6]), .Y(n3651) );
  AOI22 U4235 ( .A0(disp1_sel[7]), .A1(disp1_bit7[6]), .B0(disp1_sel[0]), .B1(
        disp1_bit0[6]), .Y(n3650) );
  NAND4 U4236 ( .A(n3654), .B(n3655), .C(n3656), .D(n3657), .Y(disp1_seg[5])
         );
  AOI22 U4237 ( .A0(disp1_sel[6]), .A1(disp1_bit6[5]), .B0(disp1_sel[5]), .B1(
        disp1_bit5[5]), .Y(n3657) );
  AOI22 U4238 ( .A0(disp1_sel[4]), .A1(disp1_bit4[5]), .B0(disp1_sel[3]), .B1(
        disp1_bit3[5]), .Y(n3656) );
  AOI22 U4239 ( .A0(disp1_sel[2]), .A1(disp1_bit2[5]), .B0(disp1_sel[1]), .B1(
        disp1_bit1[5]), .Y(n3655) );
  AOI22 U4240 ( .A0(disp1_sel[7]), .A1(disp1_bit7[5]), .B0(disp1_sel[0]), .B1(
        disp1_bit0[5]), .Y(n3654) );
  NAND4 U4241 ( .A(n3658), .B(n3659), .C(n3660), .D(n3661), .Y(disp1_seg[4])
         );
  AOI22 U4242 ( .A0(disp1_sel[6]), .A1(disp1_bit6[4]), .B0(disp1_sel[5]), .B1(
        disp1_bit5[4]), .Y(n3661) );
  AOI22 U4243 ( .A0(disp1_sel[4]), .A1(disp1_bit4[4]), .B0(disp1_sel[3]), .B1(
        disp1_bit3[4]), .Y(n3660) );
  AOI22 U4244 ( .A0(disp1_sel[2]), .A1(disp1_bit2[4]), .B0(disp1_sel[1]), .B1(
        disp1_bit1[4]), .Y(n3659) );
  AOI22 U4245 ( .A0(disp1_sel[7]), .A1(disp1_bit7[4]), .B0(disp1_sel[0]), .B1(
        disp1_bit0[4]), .Y(n3658) );
  NAND4 U4246 ( .A(n3662), .B(n3663), .C(n3664), .D(n3665), .Y(disp1_seg[3])
         );
  AOI22 U4247 ( .A0(disp1_sel[6]), .A1(disp1_bit6[3]), .B0(disp1_sel[5]), .B1(
        disp1_bit5[3]), .Y(n3665) );
  AOI22 U4248 ( .A0(disp1_sel[4]), .A1(disp1_bit4[3]), .B0(disp1_sel[3]), .B1(
        disp1_bit3[3]), .Y(n3664) );
  AOI22 U4249 ( .A0(disp1_sel[2]), .A1(disp1_bit2[3]), .B0(disp1_sel[1]), .B1(
        disp1_bit1[3]), .Y(n3663) );
  AOI22 U4250 ( .A0(disp1_sel[7]), .A1(disp1_bit7[3]), .B0(disp1_sel[0]), .B1(
        disp1_bit0[3]), .Y(n3662) );
  NAND4 U4251 ( .A(n3666), .B(n3667), .C(n3668), .D(n3669), .Y(disp1_seg[2])
         );
  AOI22 U4252 ( .A0(disp1_sel[6]), .A1(disp1_bit6[2]), .B0(disp1_sel[5]), .B1(
        disp1_bit5[2]), .Y(n3669) );
  AOI22 U4253 ( .A0(disp1_sel[4]), .A1(disp1_bit4[2]), .B0(disp1_sel[3]), .B1(
        disp1_bit3[2]), .Y(n3668) );
  AOI22 U4254 ( .A0(disp1_sel[2]), .A1(disp1_bit2[2]), .B0(disp1_sel[1]), .B1(
        disp1_bit1[2]), .Y(n3667) );
  AOI22 U4255 ( .A0(disp1_sel[7]), .A1(disp1_bit7[2]), .B0(disp1_sel[0]), .B1(
        disp1_bit0[2]), .Y(n3666) );
  NAND4 U4256 ( .A(n3670), .B(n3671), .C(n3672), .D(n3673), .Y(disp1_seg[1])
         );
  AOI22 U4257 ( .A0(disp1_sel[6]), .A1(disp1_bit6[1]), .B0(disp1_sel[5]), .B1(
        disp1_bit5[1]), .Y(n3673) );
  AOI22 U4258 ( .A0(disp1_sel[4]), .A1(disp1_bit4[1]), .B0(disp1_sel[3]), .B1(
        disp1_bit3[1]), .Y(n3672) );
  AOI22 U4259 ( .A0(disp1_sel[2]), .A1(disp1_bit2[1]), .B0(disp1_sel[1]), .B1(
        disp1_bit1[1]), .Y(n3671) );
  AOI22 U4260 ( .A0(disp1_sel[7]), .A1(disp1_bit7[1]), .B0(disp1_sel[0]), .B1(
        disp1_bit0[1]), .Y(n3670) );
  NAND4 U4261 ( .A(n3674), .B(n3675), .C(n3676), .D(n3677), .Y(disp1_seg[0])
         );
  AOI22 U4262 ( .A0(disp1_sel[6]), .A1(disp1_bit6[0]), .B0(disp1_sel[5]), .B1(
        disp1_bit5[0]), .Y(n3677) );
  NOR2B U4263 ( .AN(n3678), .B(n4978), .Y(n4990) );
  NOR2B U4264 ( .AN(n3679), .B(n3680), .Y(n4989) );
  AOI22 U4265 ( .A0(disp1_sel[4]), .A1(disp1_bit4[0]), .B0(disp1_sel[3]), .B1(
        disp1_bit3[0]), .Y(n3676) );
  NOR2B U4266 ( .AN(n3678), .B(disp1_sel_cnt[0]), .Y(n4991) );
  AOI22 U4267 ( .A0(disp1_sel[2]), .A1(disp1_bit2[0]), .B0(disp1_sel[1]), .B1(
        disp1_bit1[0]), .Y(n3675) );
  NOR2B U4268 ( .AN(n3681), .B(n4978), .Y(n4994) );
  NOR2B U4269 ( .AN(n3679), .B(disp1_sel_cnt[2]), .Y(n4993) );
  AOI22 U4270 ( .A0(disp1_sel[7]), .A1(disp1_bit7[0]), .B0(disp1_sel[0]), .B1(
        disp1_bit0[0]), .Y(n3674) );
  NOR2B U4271 ( .AN(n3429), .B(out_sel_cnt[0]), .Y(N5398) );
  NOR2 U4272 ( .A(out_sel_cnt[2]), .B(out_sel_cnt[1]), .Y(n3429) );
  NOR2B U4273 ( .AN(n3649), .B(disp2_sel_cnt[0]), .Y(N5346) );
  NOR2 U4274 ( .A(disp2_sel_cnt[1]), .B(disp2_sel_cnt[2]), .Y(n3649) );
  NOR3B U4275 ( .AN(disp2_sel_cnt[1]), .B(n4979), .C(n3648), .Y(N5323) );
  OAI211 U4276 ( .A0(disp2_sel_cnt[0]), .A1(n3648), .B0(n2728), .C0(n3682), 
        .Y(N5321) );
  INV U4277 ( .A(n3646), .Y(n3682) );
  NOR2 U4278 ( .A(disp2_sel_cnt[1]), .B(n3648), .Y(n3646) );
  NOR3B U4279 ( .AN(disp2_sel_cnt[1]), .B(disp2_sel_cnt[2]), .C(n4979), .Y(
        n4998) );
  INV U4280 ( .A(disp2_sel_cnt[2]), .Y(n3648) );
  OAI21 U4281 ( .A0(disp2_sel_cnt[1]), .A1(n4979), .B0(n3683), .Y(N5320) );
  INV U4282 ( .A(n3647), .Y(n3683) );
  NOR2B U4283 ( .AN(disp2_sel_cnt[1]), .B(disp2_sel_cnt[0]), .Y(n3647) );
  INV U4284 ( .A(disp2_sel_cnt[0]), .Y(n4979) );
  NOR2B U4285 ( .AN(n3681), .B(disp1_sel_cnt[0]), .Y(N5294) );
  NOR2 U4286 ( .A(disp1_sel_cnt[1]), .B(disp1_sel_cnt[2]), .Y(n3681) );
  NOR3B U4287 ( .AN(disp1_sel_cnt[1]), .B(n4978), .C(n3680), .Y(N5271) );
  OAI211 U4288 ( .A0(disp1_sel_cnt[0]), .A1(n3680), .B0(n2722), .C0(n3684), 
        .Y(N5269) );
  INV U4289 ( .A(n3678), .Y(n3684) );
  NOR2 U4290 ( .A(disp1_sel_cnt[1]), .B(n3680), .Y(n3678) );
  NOR3B U4291 ( .AN(disp1_sel_cnt[1]), .B(disp1_sel_cnt[2]), .C(n4978), .Y(
        n4992) );
  INV U4292 ( .A(disp1_sel_cnt[2]), .Y(n3680) );
  OAI21 U4293 ( .A0(disp1_sel_cnt[1]), .A1(n4978), .B0(n3685), .Y(N5268) );
  INV U4294 ( .A(n3679), .Y(n3685) );
  NOR2B U4295 ( .AN(disp1_sel_cnt[1]), .B(disp1_sel_cnt[0]), .Y(n3679) );
  INV U4296 ( .A(disp1_sel_cnt[0]), .Y(n4978) );
  INV U4297 ( .A(n3686), .Y(N5264) );
  NOR4B U4298 ( .AN(n3687), .B(n3688), .C(n3689), .D(n3690), .Y(n3686) );
  MX2 U4299 ( .A(n3691), .B(n3692), .S0(n3693), .Y(n3690) );
  OAI21 U4300 ( .A0(n2647), .A1(n3695), .B0(n2691), .Y(n3692) );
  OAI222 U4301 ( .A0(n2646), .A1(n3697), .B0(n3698), .B1(n2691), .C0(n3699), 
        .C1(n3700), .Y(n3689) );
  NOR2B U4302 ( .AN(n3701), .B(n3702), .Y(n3699) );
  MX2 U4303 ( .A(n3703), .B(n3704), .S0(n3705), .Y(n3688) );
  OAI21 U4304 ( .A0(n3702), .A1(n3706), .B0(n2684), .Y(n3704) );
  NOR2B U4305 ( .AN(n2684), .B(n3707), .Y(n3703) );
  OAI211 U4306 ( .A0(n3708), .A1(n3709), .B0(n3687), .C0(n3710), .Y(N5263) );
  INV U4307 ( .A(n3711), .Y(n3710) );
  OAI222 U4308 ( .A0(n3712), .A1(n3695), .B0(n3698), .B1(n3713), .C0(n3701), 
        .C1(n3714), .Y(n3711) );
  NOR2 U4309 ( .A(n3715), .B(n3707), .Y(n3714) );
  NOR2B U4310 ( .AN(n3716), .B(n3717), .Y(n3713) );
  INV U4311 ( .A(n3691), .Y(n3712) );
  INV U4312 ( .A(n3718), .Y(n3709) );
  INV U4313 ( .A(n3719), .Y(N5262) );
  NOR4B U4314 ( .AN(n3720), .B(n3718), .C(n3721), .D(n3722), .Y(n3719) );
  OAI22 U4315 ( .A0(n3723), .A1(n3701), .B0(n3724), .B1(n3695), .Y(n3722) );
  OAI2BB2 U4316 ( .B0(n3725), .B1(n3698), .A0N(n2684), .A1N(n3708), .Y(n3721)
         );
  OAI211 U4317 ( .A0(n3697), .A1(n3726), .B0(n3727), .C0(n3728), .Y(N5261) );
  NOR4 U4318 ( .A(n3691), .B(n3729), .C(n3730), .D(n3731), .Y(n3728) );
  MX2 U4319 ( .A(n3732), .B(n3733), .S0(data_type), .Y(n3731) );
  NOR2B U4320 ( .AN(n3715), .B(n3702), .Y(n3733) );
  AOI2BB1 U4321 ( .A0N(n2684), .A1N(n3700), .B0(n3718), .Y(n3715) );
  NOR2 U4322 ( .A(n3693), .B(n3716), .Y(n3732) );
  XOR2 U4323 ( .A(n2691), .B(n3695), .Y(n3716) );
  AOI2BB1 U4324 ( .A0N(n3700), .A1N(n3734), .B0(n3708), .Y(n3730) );
  NOR2 U4325 ( .A(n2684), .B(n3707), .Y(n3734) );
  NOR3 U4326 ( .A(n2684), .B(n3700), .C(n3701), .Y(n3729) );
  NOR2B U4327 ( .AN(n2647), .B(n2690), .Y(n3691) );
  NOR2 U4328 ( .A(n3735), .B(n3736), .Y(n3726) );
  NOR2B U4329 ( .AN(n2647), .B(n3717), .Y(n3736) );
  NOR2 U4330 ( .A(n2691), .B(n3698), .Y(n3735) );
  OAI211 U4331 ( .A0(n3707), .A1(n3708), .B0(n3687), .C0(n3737), .Y(N5260) );
  NOR2B U4332 ( .AN(n3738), .B(n3739), .Y(n3737) );
  AOI222 U4333 ( .A0(n3706), .A1(n3740), .B0(n2647), .B1(n3693), .C0(n2690), 
        .C1(n3741), .Y(n3738) );
  AOI22 U4334 ( .A0(n3741), .A1(n3717), .B0(n3740), .B1(n3707), .Y(n3687) );
  INV U4335 ( .A(n3742), .Y(N5259) );
  NOR4BB U4336 ( .AN(n3720), .BN(n3743), .C(n3744), .D(n3739), .Y(n3742) );
  NOR2B U4337 ( .AN(n3740), .B(n3723), .Y(n3744) );
  NOR2 U4338 ( .A(n2684), .B(n4961), .Y(n3740) );
  AOI222 U4339 ( .A0(n3745), .A1(n3741), .B0(n2691), .B1(n3746), .C0(n3700), 
        .C1(n3747), .Y(n3743) );
  NOR2 U4340 ( .A(n3707), .B(n3701), .Y(n3747) );
  NOR2 U4341 ( .A(n3698), .B(n3717), .Y(n3746) );
  NOR2 U4342 ( .A(data_type), .B(n3697), .Y(n3741) );
  INV U4343 ( .A(n3725), .Y(n3745) );
  NAND2 U4344 ( .A(n3727), .B(n3748), .Y(N5258) );
  NOR4BB U4345 ( .AN(n3720), .BN(n3749), .C(n3739), .D(n3750), .Y(n3748) );
  OAI33 U4346 ( .A0(n3707), .A1(n2684), .A2(n3701), .B0(n3717), .B1(n3697), 
        .B2(n3698), .Y(n3750) );
  OR2 U4347 ( .A(data_type), .B(n2647), .Y(n3698) );
  INV U4348 ( .A(n3695), .Y(n3697) );
  NAND2B U4349 ( .AN(n3705), .B(data_type), .Y(n3701) );
  OAI21 U4350 ( .A0(n3700), .A1(n3708), .B0(n3751), .Y(n3739) );
  INV U4351 ( .A(n3724), .Y(n3751) );
  NOR2B U4352 ( .AN(n2647), .B(n2691), .Y(n3724) );
  INV U4353 ( .A(n3705), .Y(n3708) );
  NOR2 U4354 ( .A(n3725), .B(n3723), .Y(n3749) );
  NOR2 U4355 ( .A(n3702), .B(n3700), .Y(n3723) );
  INV U4356 ( .A(n3706), .Y(n3700) );
  NOR2 U4357 ( .A(n2691), .B(n3693), .Y(n3725) );
  INV U4358 ( .A(n3717), .Y(n3693) );
  AOI22 U4359 ( .A0(n2647), .A1(n3717), .B0(n3705), .B1(n3707), .Y(n3720) );
  NOR2 U4360 ( .A(n3752), .B(n2734), .Y(n3705) );
  NOR2B U4361 ( .AN(n2721), .B(n3752), .Y(n3694) );
  NOR2 U4362 ( .A(\uut/mant_out[3] ), .B(error), .Y(n3752) );
  AOI22 U4363 ( .A0(n3702), .A1(n3718), .B0(n2691), .B1(n3753), .Y(n3727) );
  NOR2 U4364 ( .A(n3695), .B(n3717), .Y(n3753) );
  NAND2B U4365 ( .AN(n3754), .B(n2721), .Y(n3717) );
  NAND2B U4366 ( .AN(n3755), .B(n2721), .Y(n3695) );
  AOI21 U4367 ( .A0(n2721), .A1(\uut/mant_out[1] ), .B0(n3756), .Y(n3696) );
  NOR2B U4368 ( .AN(n2684), .B(n3706), .Y(n3718) );
  OAI21 U4369 ( .A0(n2734), .A1(n3609), .B0(n2747), .Y(n3706) );
  INV U4370 ( .A(\uut/mant_out[1] ), .Y(n3609) );
  NOR2 U4371 ( .A(\uut/mant_out[0] ), .B(error), .Y(n3755) );
  INV U4372 ( .A(n3707), .Y(n3702) );
  NAND2B U4373 ( .AN(n3754), .B(n2735), .Y(n3707) );
  NOR2 U4374 ( .A(\uut/mant_out[2] ), .B(error), .Y(n3754) );
  INV U4375 ( .A(n3758), .Y(N5150) );
  NOR4B U4376 ( .AN(n3759), .B(n3760), .C(n3761), .D(n3762), .Y(n3758) );
  MX2 U4377 ( .A(n3763), .B(n3764), .S0(n3765), .Y(n3762) );
  OAI21 U4378 ( .A0(n2649), .A1(n3767), .B0(n2693), .Y(n3764) );
  OAI222 U4379 ( .A0(n2648), .A1(n3769), .B0(n3770), .B1(n2693), .C0(n3771), 
        .C1(n3772), .Y(n3761) );
  NOR2B U4380 ( .AN(n3773), .B(n3774), .Y(n3771) );
  MX2 U4381 ( .A(n3775), .B(n3776), .S0(n3777), .Y(n3760) );
  OAI21 U4382 ( .A0(n3774), .A1(n3778), .B0(n2685), .Y(n3776) );
  NOR2B U4383 ( .AN(n2685), .B(n3779), .Y(n3775) );
  OAI211 U4384 ( .A0(n3780), .A1(n3781), .B0(n3759), .C0(n3782), .Y(N5149) );
  INV U4385 ( .A(n3783), .Y(n3782) );
  OAI222 U4386 ( .A0(n3784), .A1(n3767), .B0(n3770), .B1(n3785), .C0(n3773), 
        .C1(n3786), .Y(n3783) );
  NOR2 U4387 ( .A(n3787), .B(n3779), .Y(n3786) );
  NOR2B U4388 ( .AN(n3788), .B(n3789), .Y(n3785) );
  INV U4389 ( .A(n3763), .Y(n3784) );
  INV U4390 ( .A(n3790), .Y(n3781) );
  INV U4391 ( .A(n3791), .Y(N5148) );
  NOR4B U4392 ( .AN(n3792), .B(n3790), .C(n3793), .D(n3794), .Y(n3791) );
  OAI22 U4393 ( .A0(n3795), .A1(n3773), .B0(n3796), .B1(n3767), .Y(n3794) );
  OAI2BB2 U4394 ( .B0(n3797), .B1(n3770), .A0N(n2685), .A1N(n3780), .Y(n3793)
         );
  OAI211 U4395 ( .A0(n3769), .A1(n3798), .B0(n3799), .C0(n3800), .Y(N5147) );
  NOR4 U4396 ( .A(n3763), .B(n3801), .C(n3802), .D(n3803), .Y(n3800) );
  MX2 U4397 ( .A(n3804), .B(n3805), .S0(data_type), .Y(n3803) );
  NOR2B U4398 ( .AN(n3787), .B(n3774), .Y(n3805) );
  AOI2BB1 U4399 ( .A0N(n2685), .A1N(n3772), .B0(n3790), .Y(n3787) );
  NOR2 U4400 ( .A(n3765), .B(n3788), .Y(n3804) );
  XOR2 U4401 ( .A(n2693), .B(n3767), .Y(n3788) );
  AOI2BB1 U4402 ( .A0N(n3772), .A1N(n3806), .B0(n3780), .Y(n3802) );
  NOR2 U4403 ( .A(n2685), .B(n3779), .Y(n3806) );
  NOR3 U4404 ( .A(n2685), .B(n3772), .C(n3773), .Y(n3801) );
  NOR2B U4405 ( .AN(n2649), .B(n2692), .Y(n3763) );
  NOR2 U4406 ( .A(n3807), .B(n3808), .Y(n3798) );
  NOR2B U4407 ( .AN(n2649), .B(n3789), .Y(n3808) );
  NOR2 U4408 ( .A(n2693), .B(n3770), .Y(n3807) );
  OAI211 U4409 ( .A0(n3779), .A1(n3780), .B0(n3759), .C0(n3809), .Y(N5146) );
  NOR2B U4410 ( .AN(n3810), .B(n3811), .Y(n3809) );
  AOI222 U4411 ( .A0(n3778), .A1(n3812), .B0(n2649), .B1(n3765), .C0(n2692), 
        .C1(n3813), .Y(n3810) );
  AOI22 U4412 ( .A0(n3813), .A1(n3789), .B0(n3812), .B1(n3779), .Y(n3759) );
  INV U4413 ( .A(n3814), .Y(N5145) );
  NOR4BB U4414 ( .AN(n3792), .BN(n3815), .C(n3816), .D(n3811), .Y(n3814) );
  NOR2B U4415 ( .AN(n3812), .B(n3795), .Y(n3816) );
  NOR2 U4416 ( .A(n2685), .B(n4961), .Y(n3812) );
  AOI222 U4417 ( .A0(n3817), .A1(n3813), .B0(n2693), .B1(n3818), .C0(n3772), 
        .C1(n3819), .Y(n3815) );
  NOR2 U4418 ( .A(n3779), .B(n3773), .Y(n3819) );
  NOR2 U4419 ( .A(n3770), .B(n3789), .Y(n3818) );
  NOR2 U4420 ( .A(data_type), .B(n3769), .Y(n3813) );
  INV U4421 ( .A(n3797), .Y(n3817) );
  NAND2 U4422 ( .A(n3799), .B(n3820), .Y(N5144) );
  NOR4BB U4423 ( .AN(n3792), .BN(n3821), .C(n3811), .D(n3822), .Y(n3820) );
  OAI33 U4424 ( .A0(n3779), .A1(n2685), .A2(n3773), .B0(n3789), .B1(n3769), 
        .B2(n3770), .Y(n3822) );
  OR2 U4425 ( .A(data_type), .B(n2649), .Y(n3770) );
  INV U4426 ( .A(n3767), .Y(n3769) );
  NAND2B U4427 ( .AN(n3777), .B(data_type), .Y(n3773) );
  OAI21 U4428 ( .A0(n3772), .A1(n3780), .B0(n3823), .Y(n3811) );
  INV U4429 ( .A(n3796), .Y(n3823) );
  NOR2B U4430 ( .AN(n2649), .B(n2693), .Y(n3796) );
  INV U4431 ( .A(n3777), .Y(n3780) );
  NOR2 U4432 ( .A(n3797), .B(n3795), .Y(n3821) );
  NOR2 U4433 ( .A(n3774), .B(n3772), .Y(n3795) );
  INV U4434 ( .A(n3778), .Y(n3772) );
  NOR2 U4435 ( .A(n2693), .B(n3765), .Y(n3797) );
  INV U4436 ( .A(n3789), .Y(n3765) );
  AOI22 U4437 ( .A0(n2649), .A1(n3789), .B0(n3777), .B1(n3779), .Y(n3792) );
  NOR2 U4438 ( .A(n3824), .B(n2734), .Y(n3777) );
  NOR2B U4439 ( .AN(n2721), .B(n3824), .Y(n3766) );
  NOR2 U4440 ( .A(\uut/mant_out[7] ), .B(error), .Y(n3824) );
  AOI22 U4441 ( .A0(n3774), .A1(n3790), .B0(n2693), .B1(n3825), .Y(n3799) );
  NOR2 U4442 ( .A(n3767), .B(n3789), .Y(n3825) );
  NAND2B U4443 ( .AN(n3826), .B(n2721), .Y(n3789) );
  NAND2B U4444 ( .AN(n3827), .B(n2721), .Y(n3767) );
  AOI21 U4445 ( .A0(n2721), .A1(\uut/mant_out[5] ), .B0(n3756), .Y(n3768) );
  NOR2B U4446 ( .AN(n2685), .B(n3778), .Y(n3790) );
  OAI21 U4447 ( .A0(n2734), .A1(n3613), .B0(n2747), .Y(n3778) );
  INV U4448 ( .A(\uut/mant_out[5] ), .Y(n3613) );
  NOR2 U4449 ( .A(\uut/mant_out[4] ), .B(error), .Y(n3827) );
  INV U4450 ( .A(n3779), .Y(n3774) );
  NAND2B U4451 ( .AN(n3826), .B(n2735), .Y(n3779) );
  NOR2 U4452 ( .A(\uut/mant_out[6] ), .B(error), .Y(n3826) );
  INV U4453 ( .A(n3828), .Y(N5036) );
  NOR4B U4454 ( .AN(n3829), .B(n3830), .C(n3831), .D(n3832), .Y(n3828) );
  OAI22 U4455 ( .A0(n2695), .A1(n3834), .B0(n3835), .B1(n2715), .Y(n3832) );
  AOI21 U4456 ( .A0(n2720), .A1(n2715), .B0(n3838), .Y(n3834) );
  NOR2 U4457 ( .A(n2720), .B(n3839), .Y(n3831) );
  NOR2B U4458 ( .AN(n2715), .B(n3840), .Y(n3839) );
  AOI211 U4459 ( .A0(n2701), .A1(n3842), .B0(n3843), .C0(n3844), .Y(n3829) );
  MX2 U4460 ( .A(n3845), .B(n3846), .S0(n2639), .Y(n3844) );
  OAI21 U4461 ( .A0(n2701), .A1(n3842), .B0(n3848), .Y(n3845) );
  INV U4462 ( .A(n3849), .Y(N5035) );
  AOI211 U4463 ( .A0(n3850), .A1(n2694), .B0(n3843), .C0(n3851), .Y(n3849) );
  OAI222 U4464 ( .A0(n3835), .A1(n3852), .B0(n3853), .B1(n3854), .C0(n3855), 
        .C1(n2701), .Y(n3851) );
  NOR2 U4465 ( .A(n3830), .B(n3846), .Y(n3855) );
  AOI21 U4466 ( .A0(n3848), .A1(n2701), .B0(n2639), .Y(n3854) );
  INV U4467 ( .A(n3856), .Y(n3853) );
  NOR2 U4468 ( .A(n2720), .B(n3857), .Y(n3852) );
  OAI211 U4469 ( .A0(n3858), .A1(n3835), .B0(n3859), .C0(n3860), .Y(N5034) );
  AOI211 U4470 ( .A0(n3856), .A1(n3861), .B0(n3840), .C0(n3862), .Y(n3860) );
  NOR2B U4471 ( .AN(n2695), .B(n3838), .Y(n3840) );
  AOI2BB1 U4472 ( .A0N(n2701), .A1N(n3863), .B0(n3850), .Y(n3859) );
  INV U4473 ( .A(n3864), .Y(N5033) );
  NOR4B U4474 ( .AN(n3865), .B(n3866), .C(n3867), .D(n3868), .Y(n3864) );
  MX2 U4475 ( .A(n3869), .B(n3870), .S0(n2695), .Y(n3868) );
  OAI2BB1 U4476 ( .A0N(n3838), .A1N(n2719), .B0(n2714), .Y(n3869) );
  OAI31 U4477 ( .A0(n3871), .A1(n2638), .A2(n3872), .B0(n3873), .Y(n3866) );
  AOI31 U4478 ( .A0(n2720), .A1(n3857), .A2(n4961), .B0(n3846), .Y(n3873) );
  NOR2 U4479 ( .A(n3874), .B(n3871), .Y(n3846) );
  XNOR2 U4480 ( .A(n3838), .B(n2715), .Y(n3857) );
  MX2 U4481 ( .A(n3861), .B(n3875), .S0(n2701), .Y(n3865) );
  NOR2 U4482 ( .A(n3830), .B(n3876), .Y(n3875) );
  NOR2B U4483 ( .AN(n3856), .B(n3848), .Y(n3830) );
  INV U4484 ( .A(n3877), .Y(N5032) );
  NOR4BB U4485 ( .AN(n3878), .BN(n3879), .C(n3880), .D(n3843), .Y(n3877) );
  OAI2BB2 U4486 ( .B0(n2638), .B1(n3872), .A0N(n2720), .A1N(n3881), .Y(n3843)
         );
  NOR2 U4487 ( .A(n2720), .B(n2695), .Y(n3880) );
  AOI211 U4488 ( .A0(n3882), .A1(n3871), .B0(n3870), .C0(n3876), .Y(n3878) );
  NOR2 U4489 ( .A(n3874), .B(n2639), .Y(n3876) );
  NOR2B U4490 ( .AN(n3881), .B(n2715), .Y(n3870) );
  INV U4491 ( .A(n3872), .Y(n3882) );
  OAI211 U4492 ( .A0(n3883), .A1(n3872), .B0(n3884), .C0(n3885), .Y(N5031) );
  AOI222 U4493 ( .A0(n3886), .A1(n3881), .B0(n3887), .B1(n3888), .C0(n3856), 
        .C1(n3889), .Y(n3884) );
  NOR2 U4494 ( .A(n2639), .B(n3871), .Y(n3889) );
  NOR2B U4495 ( .AN(n2715), .B(n2720), .Y(n3888) );
  INV U4496 ( .A(n3835), .Y(n3887) );
  NAND2B U4497 ( .AN(data_type), .B(n2695), .Y(n3835) );
  INV U4498 ( .A(n3858), .Y(n3886) );
  NAND2 U4499 ( .A(data_type), .B(n2701), .Y(n3872) );
  NAND3 U4500 ( .A(n3885), .B(n3890), .C(n3891), .Y(N5030) );
  AOI211 U4501 ( .A0(n3881), .A1(n3892), .B0(n3883), .C0(n3858), .Y(n3891) );
  NOR2B U4502 ( .AN(n2720), .B(n2715), .Y(n3858) );
  INV U4503 ( .A(n3861), .Y(n3883) );
  NAND2 U4504 ( .A(n2639), .B(n3871), .Y(n3861) );
  INV U4505 ( .A(n3848), .Y(n3871) );
  NOR2B U4506 ( .AN(n2695), .B(n2720), .Y(n3892) );
  NOR2B U4507 ( .AN(n3838), .B(data_type), .Y(n3881) );
  AOI31 U4508 ( .A0(n3856), .A1(n2701), .A2(n2638), .B0(n3867), .Y(n3890) );
  OAI2BB2 U4509 ( .B0(n2720), .B1(n3893), .A0N(n3848), .A1N(n3894), .Y(n3867)
         );
  NOR2 U4510 ( .A(n2639), .B(n2701), .Y(n3894) );
  INV U4511 ( .A(n3850), .Y(n3893) );
  NOR2B U4512 ( .AN(n2715), .B(n3838), .Y(n3850) );
  AOI21 U4513 ( .A0(\uut/mant_out[8] ), .A1(n2547), .B0(n3756), .Y(n3838) );
  NOR2B U4514 ( .AN(n2721), .B(n2736), .Y(n3756) );
  AOI21 U4515 ( .A0(n2735), .A1(\uut/mant_out[8] ), .B0(n2748), .Y(n3841) );
  NOR2 U4516 ( .A(n4961), .B(n3842), .Y(n3856) );
  INV U4517 ( .A(n3874), .Y(n3842) );
  NOR2B U4518 ( .AN(n3879), .B(n3862), .Y(n3885) );
  OAI22 U4519 ( .A0(n3874), .A1(n2638), .B0(n2695), .B1(n2719), .Y(n3862) );
  AOI21 U4520 ( .A0(n2547), .A1(\uut/exp_out[0] ), .B0(n3897), .Y(n3837) );
  AOI21 U4521 ( .A0(n2735), .A1(\uut/mant_out[10] ), .B0(n2748), .Y(n3847) );
  AOI2BB1 U4522 ( .A0N(n2695), .A1N(n2715), .B0(n3863), .Y(n3879) );
  NOR2 U4523 ( .A(n3848), .B(n3874), .Y(n3863) );
  AOI21 U4524 ( .A0(n2735), .A1(\uut/mant_out[11] ), .B0(n2748), .Y(n3874) );
  AOI21 U4525 ( .A0(n2735), .A1(\uut/mant_out[9] ), .B0(n2748), .Y(n3848) );
  OAI21 U4526 ( .A0(\uut/mant_out[9] ), .A1(error), .B0(n2721), .Y(n3836) );
  AOI21 U4527 ( .A0(n2547), .A1(\uut/exp_out[1] ), .B0(n3897), .Y(n3833) );
  OR4 U4528 ( .A(n3898), .B(n3899), .C(n3900), .D(n3901), .Y(N4922) );
  MX2 U4529 ( .A(n3902), .B(n3903), .S0(n3904), .Y(n3901) );
  OAI21 U4530 ( .A0(n3905), .A1(n2687), .B0(n2665), .Y(n3903) );
  NOR2B U4531 ( .AN(n2665), .B(n3908), .Y(n3902) );
  MX2 U4532 ( .A(n3909), .B(n3910), .S0(n3911), .Y(n3900) );
  OAI2BB1 U4533 ( .A0N(n2552), .A1N(n2689), .B0(n2550), .Y(n3910) );
  NOR2 U4534 ( .A(n2552), .B(n2551), .Y(n3909) );
  OAI22 U4535 ( .A0(n3914), .A1(n2686), .B0(n2689), .B1(n3915), .Y(n3899) );
  NOR2 U4536 ( .A(n3916), .B(n2553), .Y(n3915) );
  NOR2 U4537 ( .A(n3905), .B(n3918), .Y(n3914) );
  INV U4538 ( .A(n3919), .Y(N4921) );
  AOI211 U4539 ( .A0(n3920), .A1(n3904), .B0(n3898), .C0(n3921), .Y(n3919) );
  OAI222 U4540 ( .A0(n3922), .A1(n3923), .B0(n3924), .B1(n3925), .C0(n3926), 
        .C1(n3927), .Y(n3921) );
  NOR2 U4541 ( .A(n2552), .B(n3928), .Y(n3927) );
  NOR2 U4542 ( .A(n3929), .B(n3908), .Y(n3925) );
  INV U4543 ( .A(n3930), .Y(n3922) );
  INV U4544 ( .A(n3931), .Y(N4920) );
  NOR4B U4545 ( .AN(n3932), .B(n3920), .C(n3930), .D(n3933), .Y(n3931) );
  OAI2BB2 U4546 ( .B0(n3934), .B1(n3926), .A0N(n3918), .A1N(n3935), .Y(n3933)
         );
  NOR2 U4547 ( .A(n3936), .B(n3937), .Y(n3932) );
  OAI2BB2 U4548 ( .B0(n2551), .B1(n3911), .A0N(n2665), .A1N(n3938), .Y(n3937)
         );
  OAI211 U4549 ( .A0(n2687), .A1(n3938), .B0(n3939), .C0(n3940), .Y(N4919) );
  NOR2 U4550 ( .A(n3941), .B(n3942), .Y(n3940) );
  OAI222 U4551 ( .A0(n3926), .A1(n3943), .B0(n2665), .B1(n3944), .C0(n3923), 
        .C1(n3945), .Y(n3942) );
  NOR2 U4552 ( .A(n2689), .B(n3946), .Y(n3945) );
  AOI21 U4553 ( .A0(n2687), .A1(n3918), .B0(n3947), .Y(n3944) );
  INV U4554 ( .A(n3948), .Y(n3943) );
  MX2 U4555 ( .A(n3949), .B(n3950), .S0(data_type), .Y(n3941) );
  NOR2B U4556 ( .AN(n3929), .B(n3905), .Y(n3950) );
  NOR2 U4557 ( .A(n3951), .B(n3920), .Y(n3929) );
  NOR2B U4558 ( .AN(n2687), .B(n2665), .Y(n3951) );
  NOR2B U4559 ( .AN(n3928), .B(n2553), .Y(n3949) );
  NOR2 U4560 ( .A(n3930), .B(n3948), .Y(n3928) );
  NOR2B U4561 ( .AN(n2551), .B(n2689), .Y(n3948) );
  OR4 U4562 ( .A(n3947), .B(n3898), .C(n3952), .D(n3953), .Y(N4918) );
  OAI222 U4563 ( .A0(n2686), .A1(n3954), .B0(n3923), .B1(n2552), .C0(n3955), 
        .C1(n2689), .Y(n3952) );
  INV U4564 ( .A(n3956), .Y(n3954) );
  OAI2BB2 U4565 ( .B0(n2553), .B1(n3955), .A0N(n3956), .A1N(n3908), .Y(n3898)
         );
  NOR2B U4566 ( .AN(n3904), .B(n3908), .Y(n3947) );
  OAI211 U4567 ( .A0(n3934), .A1(n3955), .B0(n3957), .C0(n3958), .Y(N4917) );
  AOI222 U4568 ( .A0(n3935), .A1(n3956), .B0(n3918), .B1(n3959), .C0(n3916), 
        .C1(n3960), .Y(n3957) );
  NOR2B U4569 ( .AN(n2689), .B(n2552), .Y(n3960) );
  INV U4570 ( .A(n3926), .Y(n3916) );
  NOR2 U4571 ( .A(n2687), .B(n3908), .Y(n3959) );
  NOR2 U4572 ( .A(n2665), .B(n4961), .Y(n3956) );
  NAND2B U4573 ( .AN(data_type), .B(n2551), .Y(n3955) );
  NAND2B U4574 ( .AN(n3961), .B(n3962), .Y(N4916) );
  NOR4BB U4575 ( .AN(n3939), .BN(n3935), .C(n3934), .D(n3963), .Y(n3962) );
  NOR2B U4576 ( .AN(n3946), .B(n3926), .Y(n3963) );
  OR2 U4577 ( .A(data_type), .B(n3911), .Y(n3926) );
  NOR2B U4578 ( .AN(n2551), .B(n2552), .Y(n3946) );
  NOR2 U4579 ( .A(n2689), .B(n2553), .Y(n3934) );
  NAND2 U4580 ( .A(n2687), .B(n3908), .Y(n3935) );
  AOI22 U4581 ( .A0(n3920), .A1(n3905), .B0(n3930), .B1(n2553), .Y(n3939) );
  NOR2B U4582 ( .AN(n2689), .B(n2551), .Y(n3930) );
  AOI21 U4583 ( .A0(n2547), .A1(\uut/exp_out[2] ), .B0(n3897), .Y(n3913) );
  NOR2B U4584 ( .AN(n2665), .B(n2687), .Y(n3920) );
  OAI31 U4585 ( .A0(n2665), .A1(n3908), .A2(n3924), .B0(n3958), .Y(n3961) );
  NOR2 U4586 ( .A(n3936), .B(n3953), .Y(n3958) );
  OAI2BB2 U4587 ( .B0(n2689), .B1(n3923), .A0N(n2687), .A1N(n3904), .Y(n3953)
         );
  AOI2BB1 U4588 ( .A0N(\uut/mant_out[13] ), .A1N(n2748), .B0(n3964), .Y(n3906)
         );
  AOI21 U4589 ( .A0(n2547), .A1(\uut/exp_out[3] ), .B0(n3897), .Y(n3912) );
  OAI22 U4590 ( .A0(n3905), .A1(n3938), .B0(n2553), .B1(n3923), .Y(n3936) );
  INV U4591 ( .A(n3911), .Y(n3923) );
  NOR2B U4592 ( .AN(n2547), .B(n3965), .Y(n3911) );
  OAI2BB1 U4593 ( .A0N(n2547), .A1N(\uut/exp_out[4] ), .B0(n3966), .Y(n3917)
         );
  INV U4594 ( .A(n3897), .Y(n3966) );
  NOR2 U4595 ( .A(data_type), .B(n3967), .Y(n3897) );
  NOR2B U4596 ( .AN(n2721), .B(error), .Y(n3895) );
  INV U4597 ( .A(n2789), .Y(n2788) );
  INV U4598 ( .A(n3918), .Y(n3924) );
  NOR2 U4599 ( .A(n3904), .B(n4961), .Y(n3918) );
  INV U4600 ( .A(n3938), .Y(n3904) );
  OAI21 U4601 ( .A0(\uut/mant_out[15] ), .A1(n2748), .B0(n3968), .Y(n3938) );
  INV U4602 ( .A(n3964), .Y(n3968) );
  INV U4603 ( .A(n3905), .Y(n3908) );
  AOI2BB1 U4604 ( .A0N(\uut/mant_out[14] ), .A1N(n2748), .B0(n3964), .Y(n3905)
         );
  AOI2BB1 U4605 ( .A0N(\uut/mant_out[12] ), .A1N(n2748), .B0(n3964), .Y(n3907)
         );
  NOR2 U4606 ( .A(n2748), .B(n2704), .Y(n3964) );
  OAI211 U4607 ( .A0(n2667), .A1(n3970), .B0(n3971), .C0(n3972), .Y(N4808) );
  OAI21 U4608 ( .A0(n3973), .A1(n2554), .B0(n3974), .Y(n3972) );
  NOR2 U4609 ( .A(n3975), .B(n3976), .Y(n3973) );
  MX2 U4610 ( .A(n2555), .B(n3978), .S0(n3975), .Y(n3971) );
  NOR2B U4611 ( .AN(n3979), .B(n3980), .Y(n3978) );
  OAI222 U4612 ( .A0(n3981), .A1(n3982), .B0(n3983), .B1(n3984), .C0(n3979), 
        .C1(n3976), .Y(N4807) );
  NOR2 U4613 ( .A(n3975), .B(n3985), .Y(n3984) );
  OAI222 U4614 ( .A0(n3983), .A1(n3986), .B0(n3982), .B1(n2667), .C0(n3987), 
        .C1(n3976), .Y(N4806) );
  NOR2 U4615 ( .A(n2555), .B(n2667), .Y(n3987) );
  OAI211 U4616 ( .A0(n3988), .A1(n3970), .B0(n3989), .C0(n3990), .Y(N4805) );
  AOI31 U4617 ( .A0(n3975), .A1(data_type), .A2(n3985), .B0(n3991), .Y(n3989)
         );
  INV U4618 ( .A(n3979), .Y(n3991) );
  NAND2B U4619 ( .AN(n2667), .B(n2555), .Y(n3979) );
  XNOR2 U4620 ( .A(n3976), .B(n2555), .Y(n3985) );
  AOI21 U4621 ( .A0(n3974), .A1(n2554), .B0(n3992), .Y(n3988) );
  AOI22 U4622 ( .A0(n2555), .A1(n3993), .B0(n2667), .B1(n3981), .Y(N4804) );
  NOR2 U4623 ( .A(n3994), .B(n3992), .Y(n3993) );
  NOR2 U4624 ( .A(n3975), .B(n2667), .Y(n3992) );
  NOR2B U4625 ( .AN(n3980), .B(n3982), .Y(n3994) );
  INV U4626 ( .A(n3981), .Y(n3980) );
  OAI21 U4627 ( .A0(n3986), .A1(n3981), .B0(n3995), .Y(N4803) );
  AOI21 U4628 ( .A0(n3996), .A1(n3974), .B0(n3997), .Y(n3995) );
  INV U4629 ( .A(n3983), .Y(n3974) );
  NAND2 U4630 ( .A(data_type), .B(n3976), .Y(n3981) );
  OR3 U4631 ( .A(n3986), .B(n3997), .C(n3998), .Y(N4802) );
  OAI31 U4632 ( .A0(n3975), .A1(n3970), .A2(n3983), .B0(n3990), .Y(n3998) );
  NAND2 U4633 ( .A(n3996), .B(n3970), .Y(n3990) );
  NAND2 U4634 ( .A(data_type), .B(n2667), .Y(n3983) );
  INV U4635 ( .A(n3976), .Y(n3970) );
  AOI21 U4636 ( .A0(n2735), .A1(\uut/mant_out[16] ), .B0(n2748), .Y(n3976) );
  NOR2 U4637 ( .A(n2667), .B(n3996), .Y(n3997) );
  NOR2 U4638 ( .A(n3975), .B(n2554), .Y(n3996) );
  INV U4639 ( .A(n3982), .Y(n3975) );
  AOI21 U4640 ( .A0(n2735), .A1(\uut/mant_out[19] ), .B0(n2748), .Y(n3969) );
  NOR2 U4641 ( .A(n2555), .B(n3982), .Y(n3986) );
  OAI2BB1 U4642 ( .A0N(n2735), .A1N(\uut/mant_out[18] ), .B0(n2747), .Y(n3982)
         );
  AOI21 U4643 ( .A0(n2735), .A1(\uut/mant_out[17] ), .B0(n2748), .Y(n3977) );
  OAI211 U4644 ( .A0(n2669), .A1(n4000), .B0(n4001), .C0(n4002), .Y(N4746) );
  OAI2BB1 U4645 ( .A0N(n4003), .A1N(n4004), .B0(n2542), .Y(n4002) );
  MX2 U4646 ( .A(n4005), .B(n4006), .S0(n4003), .Y(n4001) );
  NOR2B U4647 ( .AN(n4007), .B(n4008), .Y(n4006) );
  INV U4648 ( .A(n4009), .Y(n4008) );
  OR2 U4649 ( .A(n4010), .B(n4004), .Y(n4005) );
  OAI222 U4650 ( .A0(n4011), .A1(n4009), .B0(n4007), .B1(n4010), .C0(n4004), 
        .C1(n4012), .Y(N4745) );
  NOR2 U4651 ( .A(n4003), .B(n4013), .Y(n4012) );
  OAI222 U4652 ( .A0(n4011), .A1(n2669), .B0(n4004), .B1(n4014), .C0(n4015), 
        .C1(n4010), .Y(N4744) );
  NOR2 U4653 ( .A(n2669), .B(n2543), .Y(n4015) );
  OAI211 U4654 ( .A0(n4017), .A1(n4000), .B0(n4018), .C0(n4019), .Y(N4743) );
  AOI31 U4655 ( .A0(n4003), .A1(data_type), .A2(n4013), .B0(n4020), .Y(n4018)
         );
  INV U4656 ( .A(n4007), .Y(n4020) );
  NAND2B U4657 ( .AN(n2669), .B(n2543), .Y(n4007) );
  XNOR2 U4658 ( .A(n4010), .B(n2543), .Y(n4013) );
  AOI2BB2 U4659 ( .B0(n2668), .B1(n4011), .A0N(n2543), .A1N(n4004), .Y(n4017)
         );
  OAI22 U4660 ( .A0(n2669), .A1(n4021), .B0(n4022), .B1(n4009), .Y(N4742) );
  NOR2 U4661 ( .A(n4011), .B(n2542), .Y(n4021) );
  OAI21 U4662 ( .A0(n4014), .A1(n4009), .B0(n4023), .Y(N4741) );
  NOR2 U4663 ( .A(n4024), .B(n4025), .Y(n4023) );
  NOR2B U4664 ( .AN(n4022), .B(n4004), .Y(n4024) );
  NAND2 U4665 ( .A(data_type), .B(n4010), .Y(n4009) );
  OR3 U4666 ( .A(n4014), .B(n4025), .C(n4026), .Y(N4740) );
  OAI31 U4667 ( .A0(n4003), .A1(n4004), .A2(n4000), .B0(n4019), .Y(n4026) );
  NAND2 U4668 ( .A(n4022), .B(n4000), .Y(n4019) );
  INV U4669 ( .A(n4010), .Y(n4000) );
  AOI21 U4670 ( .A0(n2735), .A1(\uut/mant_out[20] ), .B0(n2748), .Y(n4010) );
  NAND2 U4671 ( .A(data_type), .B(n2669), .Y(n4004) );
  NOR2 U4672 ( .A(n2669), .B(n4022), .Y(n4025) );
  NOR2 U4673 ( .A(n4003), .B(n2542), .Y(n4022) );
  INV U4674 ( .A(n4011), .Y(n4003) );
  AOI21 U4675 ( .A0(n2704), .A1(\uut/exp_out[0] ), .B0(n4027), .Y(n3999) );
  NOR2 U4676 ( .A(n2543), .B(n4011), .Y(n4014) );
  OAI2BB1 U4677 ( .A0N(n2735), .A1N(\uut/mant_out[22] ), .B0(n2747), .Y(n4011)
         );
  AOI21 U4678 ( .A0(n2735), .A1(\uut/mant_out[21] ), .B0(n2748), .Y(n4016) );
  NOR2B U4679 ( .AN(error), .B(n2734), .Y(n3896) );
  OAI211 U4680 ( .A0(n2671), .A1(n4029), .B0(n4030), .C0(n4031), .Y(N4684) );
  OAI21 U4681 ( .A0(n4032), .A1(n2556), .B0(n4033), .Y(n4031) );
  NOR2 U4682 ( .A(n4034), .B(n4035), .Y(n4032) );
  MX2 U4683 ( .A(n2557), .B(n4037), .S0(n4034), .Y(n4030) );
  NOR2B U4684 ( .AN(n4038), .B(n4039), .Y(n4037) );
  OAI222 U4685 ( .A0(n4040), .A1(n4041), .B0(n4042), .B1(n4043), .C0(n4038), 
        .C1(n4035), .Y(N4683) );
  NOR2 U4686 ( .A(n4034), .B(n4044), .Y(n4043) );
  OAI222 U4687 ( .A0(n4042), .A1(n4045), .B0(n4041), .B1(n2671), .C0(n4046), 
        .C1(n4035), .Y(N4682) );
  NOR2 U4688 ( .A(n2557), .B(n2671), .Y(n4046) );
  OAI211 U4689 ( .A0(n4047), .A1(n4029), .B0(n4048), .C0(n4049), .Y(N4681) );
  AOI31 U4690 ( .A0(n4034), .A1(data_type), .A2(n4044), .B0(n4050), .Y(n4048)
         );
  INV U4691 ( .A(n4038), .Y(n4050) );
  NAND2B U4692 ( .AN(n2671), .B(n2557), .Y(n4038) );
  XNOR2 U4693 ( .A(n4035), .B(n2557), .Y(n4044) );
  AOI21 U4694 ( .A0(n4033), .A1(n2556), .B0(n4051), .Y(n4047) );
  AOI22 U4695 ( .A0(n2557), .A1(n4052), .B0(n2671), .B1(n4040), .Y(N4680) );
  NOR2 U4696 ( .A(n4053), .B(n4051), .Y(n4052) );
  NOR2 U4697 ( .A(n4034), .B(n2671), .Y(n4051) );
  NOR2B U4698 ( .AN(n4039), .B(n4041), .Y(n4053) );
  INV U4699 ( .A(n4040), .Y(n4039) );
  OAI21 U4700 ( .A0(n4045), .A1(n4040), .B0(n4054), .Y(N4679) );
  AOI21 U4701 ( .A0(n4055), .A1(n4033), .B0(n4056), .Y(n4054) );
  INV U4702 ( .A(n4042), .Y(n4033) );
  NAND2 U4703 ( .A(data_type), .B(n4035), .Y(n4040) );
  OR3 U4704 ( .A(n4045), .B(n4056), .C(n4057), .Y(N4678) );
  OAI31 U4705 ( .A0(n4034), .A1(n4029), .A2(n4042), .B0(n4049), .Y(n4057) );
  NAND2 U4706 ( .A(n4055), .B(n4029), .Y(n4049) );
  NAND2 U4707 ( .A(data_type), .B(n2671), .Y(n4042) );
  INV U4708 ( .A(n4035), .Y(n4029) );
  AOI21 U4709 ( .A0(n2704), .A1(\uut/exp_out[1] ), .B0(n4027), .Y(n4035) );
  NOR2 U4710 ( .A(n2671), .B(n4055), .Y(n4056) );
  NOR2 U4711 ( .A(n4034), .B(n2556), .Y(n4055) );
  INV U4712 ( .A(n4041), .Y(n4034) );
  AOI21 U4713 ( .A0(n2704), .A1(\uut/exp_out[4] ), .B0(n4027), .Y(n4028) );
  NOR2 U4714 ( .A(n2557), .B(n4041), .Y(n4045) );
  OAI2BB1 U4715 ( .A0N(n2704), .A1N(\uut/exp_out[3] ), .B0(n4058), .Y(n4041)
         );
  AOI21 U4716 ( .A0(n2704), .A1(\uut/exp_out[2] ), .B0(n4027), .Y(n4036) );
  OAI211 U4717 ( .A0(n4059), .A1(n4060), .B0(n4061), .C0(n4062), .Y(N4622) );
  OAI21 U4718 ( .A0(n4063), .A1(n2710), .B0(n4065), .Y(n4062) );
  MX2 U4719 ( .A(n4066), .B(n4067), .S0(n2710), .Y(n4061) );
  NAND2 U4720 ( .A(n4063), .B(n4060), .Y(n4067) );
  NOR2B U4721 ( .AN(n4068), .B(n4069), .Y(n4066) );
  OAI222 U4722 ( .A0(n4070), .A1(n4071), .B0(n4068), .B1(n4072), .C0(n2710), 
        .C1(n4073), .Y(N4621) );
  NOR2 U4723 ( .A(n4063), .B(n4069), .Y(n4073) );
  OAI222 U4724 ( .A0(n4059), .A1(n2710), .B0(n4072), .B1(n4074), .C0(n4070), 
        .C1(n4075), .Y(N4620) );
  NOR2B U4725 ( .AN(n4076), .B(n4077), .Y(n4074) );
  INV U4726 ( .A(n4078), .Y(N4619) );
  AOI211 U4727 ( .A0(n4072), .A1(n4079), .B0(n4080), .C0(n4081), .Y(n4078) );
  OAI31 U4728 ( .A0(n4071), .A1(n2710), .A2(n4961), .B0(n4068), .Y(n4081) );
  NAND2 U4729 ( .A(n4076), .B(n4077), .Y(n4068) );
  XNOR2 U4730 ( .A(n4072), .B(n4065), .Y(n4071) );
  OAI2BB2 U4731 ( .B0(n4077), .B1(n4070), .A0N(n4076), .A1N(n2710), .Y(n4079)
         );
  OAI22 U4732 ( .A0(n4082), .A1(n4083), .B0(n4084), .B1(n4059), .Y(N4618) );
  NOR2 U4733 ( .A(n2710), .B(n4065), .Y(n4084) );
  OAI21 U4734 ( .A0(n4075), .A1(n4083), .B0(n4085), .Y(N4617) );
  AOI21 U4735 ( .A0(n4082), .A1(n4063), .B0(n4086), .Y(n4085) );
  INV U4736 ( .A(n4070), .Y(n4063) );
  INV U4737 ( .A(n4069), .Y(n4083) );
  NOR2 U4738 ( .A(n4961), .B(n4060), .Y(n4069) );
  OR4 U4739 ( .A(n4075), .B(n4080), .C(n4086), .D(n4087), .Y(N4616) );
  NOR3B U4740 ( .AN(n2710), .B(n4070), .C(n4060), .Y(n4087) );
  INV U4741 ( .A(n4072), .Y(n4060) );
  NAND2B U4742 ( .AN(n4076), .B(data_type), .Y(n4070) );
  NOR2 U4743 ( .A(n4082), .B(n4059), .Y(n4086) );
  INV U4744 ( .A(n4076), .Y(n4059) );
  NOR2B U4745 ( .AN(n2704), .B(n3965), .Y(n4076) );
  XNOR2 U4746 ( .A(n4088), .B(n4089), .Y(n3965) );
  MX2 U4747 ( .A(\uut/in1_16_reg[15] ), .B(\uut/in1_32_reg[31] ), .S0(
        data_type), .Y(n4089) );
  MX2 U4748 ( .A(\uut/in2_16_reg[15] ), .B(\uut/in2_32_reg[31] ), .S0(
        data_type), .Y(n4088) );
  NOR2B U4749 ( .AN(n4082), .B(n4072), .Y(n4080) );
  AOI21 U4750 ( .A0(n2704), .A1(\uut/exp_out[5] ), .B0(n4027), .Y(n4072) );
  NOR2B U4751 ( .AN(n2710), .B(n4065), .Y(n4082) );
  NOR2 U4752 ( .A(n4077), .B(n2710), .Y(n4075) );
  OAI2BB1 U4753 ( .A0N(n2704), .A1N(\uut/exp_out[7] ), .B0(n4058), .Y(n4064)
         );
  INV U4754 ( .A(n4065), .Y(n4077) );
  OAI2BB1 U4755 ( .A0N(n2704), .A1N(\uut/exp_out[6] ), .B0(n4058), .Y(n4065)
         );
  INV U4756 ( .A(n4027), .Y(n4058) );
  NOR2 U4757 ( .A(n4961), .B(n3967), .Y(n4027) );
  OAI21 U4758 ( .A0(error), .A1(n4090), .B0(n4091), .Y(n3967) );
  NOR2B U4759 ( .AN(n2789), .B(n4961), .Y(n3757) );
  NOR2B U4760 ( .AN(n4091), .B(n4090), .Y(n2789) );
  OAI2BB1 U4761 ( .A0N(n3595), .A1N(n4092), .B0(n4093), .Y(n4090) );
  AOI222 U4762 ( .A0(n2537), .A1(n4094), .B0(n2535), .B1(n4096), .C0(n4097), 
        .C1(n4098), .Y(n4093) );
  INV U4763 ( .A(n3603), .Y(n4097) );
  INV U4764 ( .A(n4099), .Y(n3595) );
  AOI211 U4765 ( .A0(n2535), .A1(n3604), .B0(n4100), .C0(n4101), .Y(n4091) );
  MX2 U4766 ( .A(n4102), .B(n4103), .S0(data_type), .Y(n4101) );
  NOR2B U4767 ( .AN(n4104), .B(n4099), .Y(n4103) );
  NOR4B U4768 ( .AN(n4105), .B(\uut/in1_32_reg[24] ), .C(\uut/in1_32_reg[25] ), 
        .D(\uut/in1_32_reg[23] ), .Y(n4104) );
  NOR4B U4769 ( .AN(n4106), .B(\uut/in1_32_reg[26] ), .C(\uut/in1_32_reg[27] ), 
        .D(\uut/in1_32_reg[28] ), .Y(n4105) );
  NOR2 U4770 ( .A(\uut/in1_32_reg[29] ), .B(\uut/in1_32_reg[30] ), .Y(n4106)
         );
  NOR4B U4771 ( .AN(n4107), .B(\uut/in1_16_reg[10] ), .C(\uut/in1_16_reg[11] ), 
        .D(n2536), .Y(n4102) );
  NOR3 U4772 ( .A(\uut/in1_16_reg[14] ), .B(\uut/in1_16_reg[12] ), .C(
        \uut/in1_16_reg[13] ), .Y(n4107) );
  NOR2B U4773 ( .AN(n3602), .B(n3603), .Y(n4100) );
  NOR4BB U4774 ( .AN(n4108), .BN(n4109), .C(\uut/in2_32_reg[26] ), .D(
        \uut/in2_32_reg[27] ), .Y(n3602) );
  NOR4 U4775 ( .A(\uut/in2_32_reg[25] ), .B(\uut/in2_32_reg[24] ), .C(
        \uut/in2_32_reg[23] ), .D(n4961), .Y(n4109) );
  NOR3 U4776 ( .A(\uut/in2_32_reg[28] ), .B(\uut/in2_32_reg[29] ), .C(
        \uut/in2_32_reg[30] ), .Y(n4108) );
  NOR4B U4777 ( .AN(n4110), .B(data_type), .C(\uut/in2_16_reg[11] ), .D(
        \uut/in2_16_reg[10] ), .Y(n3604) );
  NOR3 U4778 ( .A(\uut/in2_16_reg[14] ), .B(\uut/in2_16_reg[12] ), .C(
        \uut/in2_16_reg[13] ), .Y(n4110) );
  OAI2BB1 U4779 ( .A0N(n4092), .A1N(n4099), .B0(n4111), .Y(n5007) );
  AOI222 U4780 ( .A0(n3603), .A1(n4098), .B0(n2536), .B1(n4094), .C0(n2534), 
        .C1(n4096), .Y(n4111) );
  NOR4BB U4781 ( .AN(\uut/in2_16_reg[11] ), .BN(n4112), .C(data_type), .D(
        n3585), .Y(n4096) );
  INV U4782 ( .A(\uut/in2_16_reg[10] ), .Y(n3585) );
  NOR3B U4783 ( .AN(\uut/in2_16_reg[14] ), .B(n3584), .C(n3583), .Y(n4112) );
  INV U4784 ( .A(\uut/in2_16_reg[13] ), .Y(n3583) );
  INV U4785 ( .A(\uut/in2_16_reg[12] ), .Y(n3584) );
  NOR4BB U4786 ( .AN(n4113), .BN(n4114), .C(\uut/in2_16_reg[5] ), .D(
        \uut/in2_16_reg[6] ), .Y(n4095) );
  NOR4B U4787 ( .AN(n4115), .B(\uut/in2_16_reg[2] ), .C(\uut/in2_16_reg[4] ), 
        .D(\uut/in2_16_reg[3] ), .Y(n4114) );
  NOR2 U4788 ( .A(\uut/in2_16_reg[1] ), .B(\uut/in2_16_reg[0] ), .Y(n4115) );
  NOR3 U4789 ( .A(\uut/in2_16_reg[7] ), .B(\uut/in2_16_reg[9] ), .C(
        \uut/in2_16_reg[8] ), .Y(n4113) );
  NOR4BB U4790 ( .AN(\uut/in1_16_reg[11] ), .BN(n4116), .C(data_type), .D(
        n3582), .Y(n4094) );
  INV U4791 ( .A(\uut/in1_16_reg[10] ), .Y(n3582) );
  NOR3B U4792 ( .AN(\uut/in1_16_reg[14] ), .B(n3581), .C(n3580), .Y(n4116) );
  INV U4793 ( .A(\uut/in1_16_reg[13] ), .Y(n3580) );
  INV U4794 ( .A(\uut/in1_16_reg[12] ), .Y(n3581) );
  NOR4BB U4795 ( .AN(n4117), .BN(n4118), .C(\uut/in1_16_reg[5] ), .D(
        \uut/in1_16_reg[6] ), .Y(n3594) );
  NOR4B U4796 ( .AN(n4119), .B(\uut/in1_16_reg[2] ), .C(\uut/in1_16_reg[4] ), 
        .D(\uut/in1_16_reg[3] ), .Y(n4118) );
  NOR2 U4797 ( .A(\uut/in1_16_reg[1] ), .B(\uut/in1_16_reg[0] ), .Y(n4119) );
  NOR3 U4798 ( .A(\uut/in1_16_reg[7] ), .B(\uut/in1_16_reg[9] ), .C(
        \uut/in1_16_reg[8] ), .Y(n4117) );
  NOR2B U4799 ( .AN(n4120), .B(n2802), .Y(n4098) );
  NAND2 U4800 ( .A(data_type), .B(\uut/in2_32_reg[30] ), .Y(n2802) );
  NOR4BB U4801 ( .AN(\uut/in2_32_reg[24] ), .BN(n4121), .C(n3561), .D(n3564), 
        .Y(n4120) );
  INV U4802 ( .A(\uut/in2_32_reg[23] ), .Y(n3564) );
  INV U4803 ( .A(\uut/in2_32_reg[25] ), .Y(n3561) );
  NOR4BB U4804 ( .AN(\uut/in2_32_reg[28] ), .BN(\uut/in2_32_reg[29] ), .C(
        n3559), .D(n3557), .Y(n4121) );
  INV U4805 ( .A(\uut/in2_32_reg[27] ), .Y(n3557) );
  INV U4806 ( .A(\uut/in2_32_reg[26] ), .Y(n3559) );
  NAND3 U4807 ( .A(n4122), .B(n4123), .C(n4124), .Y(n3603) );
  NOR4BB U4808 ( .AN(n4125), .BN(n4126), .C(\uut/in2_32_reg[10] ), .D(
        \uut/in2_32_reg[0] ), .Y(n4124) );
  NOR4B U4809 ( .AN(n4127), .B(\uut/in2_32_reg[17] ), .C(\uut/in2_32_reg[19] ), 
        .D(\uut/in2_32_reg[18] ), .Y(n4126) );
  NOR3 U4810 ( .A(\uut/in2_32_reg[14] ), .B(\uut/in2_32_reg[16] ), .C(
        \uut/in2_32_reg[15] ), .Y(n4127) );
  NOR3 U4811 ( .A(\uut/in2_32_reg[11] ), .B(\uut/in2_32_reg[13] ), .C(
        \uut/in2_32_reg[12] ), .Y(n4125) );
  NOR4B U4812 ( .AN(n4128), .B(\uut/in2_32_reg[22] ), .C(\uut/in2_32_reg[3] ), 
        .D(\uut/in2_32_reg[2] ), .Y(n4123) );
  NOR3 U4813 ( .A(\uut/in2_32_reg[1] ), .B(\uut/in2_32_reg[21] ), .C(
        \uut/in2_32_reg[20] ), .Y(n4128) );
  NOR4B U4814 ( .AN(n4129), .B(\uut/in2_32_reg[7] ), .C(\uut/in2_32_reg[9] ), 
        .D(\uut/in2_32_reg[8] ), .Y(n4122) );
  NOR3 U4815 ( .A(\uut/in2_32_reg[4] ), .B(\uut/in2_32_reg[6] ), .C(
        \uut/in2_32_reg[5] ), .Y(n4129) );
  NAND3 U4816 ( .A(n4130), .B(n4131), .C(n4132), .Y(n4099) );
  NOR4BB U4817 ( .AN(n4133), .BN(n4134), .C(\uut/in1_32_reg[10] ), .D(
        \uut/in1_32_reg[0] ), .Y(n4132) );
  NOR4B U4818 ( .AN(n4135), .B(\uut/in1_32_reg[17] ), .C(\uut/in1_32_reg[19] ), 
        .D(\uut/in1_32_reg[18] ), .Y(n4134) );
  NOR3 U4819 ( .A(\uut/in1_32_reg[14] ), .B(\uut/in1_32_reg[16] ), .C(
        \uut/in1_32_reg[15] ), .Y(n4135) );
  NOR3 U4820 ( .A(\uut/in1_32_reg[11] ), .B(\uut/in1_32_reg[13] ), .C(
        \uut/in1_32_reg[12] ), .Y(n4133) );
  NOR4B U4821 ( .AN(n4136), .B(\uut/in1_32_reg[22] ), .C(\uut/in1_32_reg[3] ), 
        .D(\uut/in1_32_reg[2] ), .Y(n4131) );
  NOR3 U4822 ( .A(\uut/in1_32_reg[1] ), .B(\uut/in1_32_reg[21] ), .C(
        \uut/in1_32_reg[20] ), .Y(n4136) );
  NOR4B U4823 ( .AN(n4137), .B(\uut/in1_32_reg[7] ), .C(\uut/in1_32_reg[9] ), 
        .D(\uut/in1_32_reg[8] ), .Y(n4130) );
  NOR3 U4824 ( .A(\uut/in1_32_reg[4] ), .B(\uut/in1_32_reg[6] ), .C(
        \uut/in1_32_reg[5] ), .Y(n4137) );
  NOR2B U4825 ( .AN(n4138), .B(n2803), .Y(n4092) );
  NAND2 U4826 ( .A(data_type), .B(\uut/in1_32_reg[30] ), .Y(n2803) );
  NOR4BB U4827 ( .AN(\uut/in1_32_reg[24] ), .BN(n4139), .C(n3534), .D(n3537), 
        .Y(n4138) );
  INV U4828 ( .A(\uut/in1_32_reg[23] ), .Y(n3537) );
  INV U4829 ( .A(\uut/in1_32_reg[25] ), .Y(n3534) );
  NOR4BB U4830 ( .AN(\uut/in1_32_reg[28] ), .BN(\uut/in1_32_reg[29] ), .C(
        n3532), .D(n3530), .Y(n4139) );
  INV U4831 ( .A(\uut/in1_32_reg[27] ), .Y(n3530) );
  INV U4832 ( .A(\uut/in1_32_reg[26] ), .Y(n3532) );
  OAI211 U4833 ( .A0(n2615), .A1(n4140), .B0(n4141), .C0(n4142), .Y(N4558) );
  NOR2 U4834 ( .A(n4143), .B(n4144), .Y(n4142) );
  MX2 U4835 ( .A(n4145), .B(n4146), .S0(n2617), .Y(n4144) );
  NOR2B U4836 ( .AN(in2_disp[1]), .B(n2777), .Y(n4146) );
  NOR2B U4837 ( .AN(n4147), .B(n2745), .Y(n4143) );
  NOR2 U4838 ( .A(n4148), .B(n4149), .Y(n4141) );
  NOR2B U4839 ( .AN(n4150), .B(n4151), .Y(n4149) );
  AOI21 U4840 ( .A0(n2617), .A1(n2615), .B0(in2_disp[1]), .Y(n4151) );
  OAI2BB1 U4841 ( .A0N(n2615), .A1N(n4145), .B0(n4152), .Y(N4557) );
  AOI211 U4842 ( .A0(n4153), .A1(n4154), .B0(n4148), .C0(n4155), .Y(n4152) );
  NOR2B U4843 ( .AN(n4150), .B(n4156), .Y(n4155) );
  NOR2B U4844 ( .AN(n4157), .B(n2616), .Y(n4156) );
  NOR2 U4845 ( .A(n2617), .B(n4158), .Y(n4148) );
  INV U4846 ( .A(n4159), .Y(N4556) );
  AOI211 U4847 ( .A0(n4160), .A1(n2781), .B0(n4162), .C0(n4163), .Y(n4159) );
  OAI22 U4848 ( .A0(n2617), .A1(n4140), .B0(n4164), .B1(n2746), .Y(n4163) );
  NOR2B U4849 ( .AN(n4150), .B(n4165), .Y(n4162) );
  NOR2B U4850 ( .AN(n4166), .B(n2615), .Y(n4165) );
  NOR2 U4851 ( .A(in2_disp[1]), .B(n2614), .Y(n4160) );
  OAI211 U4852 ( .A0(n2615), .A1(n4167), .B0(n4168), .C0(n4169), .Y(N4555) );
  NAND2B U4853 ( .AN(n2745), .B(n4170), .Y(n4169) );
  OAI31 U4854 ( .A0(n2677), .A1(n2604), .A2(n4171), .B0(n4172), .Y(n4170) );
  AOI211 U4855 ( .A0(n2781), .A1(n4173), .B0(n4145), .C0(n4174), .Y(n4168) );
  NOR2 U4856 ( .A(in2_disp[1]), .B(n4140), .Y(n4145) );
  NOR2 U4857 ( .A(n2617), .B(n4157), .Y(n4173) );
  XOR2 U4858 ( .A(in2_disp[1]), .B(n2615), .Y(n4157) );
  AOI22 U4859 ( .A0(n4175), .A1(n2617), .B0(n4150), .B1(in2_disp[1]), .Y(n4167) );
  OAI222 U4860 ( .A0(n4158), .A1(n4176), .B0(n2746), .B1(n4177), .C0(n4140), 
        .C1(n4178), .Y(N4554) );
  NOR2 U4861 ( .A(n2617), .B(in2_disp[1]), .Y(n4178) );
  OAI21 U4862 ( .A0(n4166), .A1(n4158), .B0(n4179), .Y(N4553) );
  AOI211 U4863 ( .A0(n4176), .A1(n4150), .B0(n4180), .C0(n4181), .Y(n4179) );
  NOR2 U4864 ( .A(n4182), .B(n2745), .Y(n4181) );
  INV U4865 ( .A(n4183), .Y(n4180) );
  NAND2B U4866 ( .AN(n2615), .B(n2781), .Y(n4158) );
  OAI211 U4867 ( .A0(n4184), .A1(n2746), .B0(n4185), .C0(n4183), .Y(N4552) );
  NAND2B U4868 ( .AN(n4176), .B(n4175), .Y(n4183) );
  INV U4869 ( .A(n4140), .Y(n4175) );
  NAND2 U4870 ( .A(in2_disp[3]), .B(n2781), .Y(n4140) );
  AOI211 U4871 ( .A0(n4150), .A1(n4186), .B0(n4174), .C0(n4187), .Y(n4185) );
  NOR2B U4872 ( .AN(n4166), .B(n2780), .Y(n4187) );
  NOR2B U4873 ( .AN(in2_disp[1]), .B(n2617), .Y(n4166) );
  NOR3B U4874 ( .AN(n4176), .B(n2778), .C(n2614), .Y(n4174) );
  NOR2B U4875 ( .AN(n2617), .B(in2_disp[1]), .Y(n4176) );
  NOR2B U4876 ( .AN(n2617), .B(n2615), .Y(n4186) );
  NOR2B U4877 ( .AN(n2781), .B(in2_disp[3]), .Y(n4150) );
  OAI211 U4878 ( .A0(n2611), .A1(n4188), .B0(n4189), .C0(n4190), .Y(N4406) );
  NOR2 U4879 ( .A(n4191), .B(n4192), .Y(n4190) );
  MX2 U4880 ( .A(n4193), .B(n4194), .S0(n2613), .Y(n4192) );
  NOR2B U4881 ( .AN(in2_disp[5]), .B(n2779), .Y(n4194) );
  NOR2B U4882 ( .AN(n4195), .B(n2745), .Y(n4191) );
  NOR2 U4883 ( .A(n4196), .B(n4197), .Y(n4189) );
  NOR2B U4884 ( .AN(n4198), .B(n4199), .Y(n4197) );
  AOI21 U4885 ( .A0(n2613), .A1(n2611), .B0(in2_disp[5]), .Y(n4199) );
  OAI2BB1 U4886 ( .A0N(n2611), .A1N(n4193), .B0(n4200), .Y(N4405) );
  AOI211 U4887 ( .A0(n4153), .A1(n4201), .B0(n4196), .C0(n4202), .Y(n4200) );
  NOR2B U4888 ( .AN(n4198), .B(n4203), .Y(n4202) );
  NOR2B U4889 ( .AN(n4204), .B(n2612), .Y(n4203) );
  NOR2 U4890 ( .A(n2613), .B(n4205), .Y(n4196) );
  INV U4891 ( .A(n4206), .Y(N4404) );
  AOI211 U4892 ( .A0(n4207), .A1(n2781), .B0(n4208), .C0(n4209), .Y(n4206) );
  OAI22 U4893 ( .A0(n2613), .A1(n4188), .B0(n4210), .B1(n2746), .Y(n4209) );
  NOR2B U4894 ( .AN(n4198), .B(n4211), .Y(n4208) );
  NOR2B U4895 ( .AN(n4212), .B(n2611), .Y(n4211) );
  NOR2 U4896 ( .A(in2_disp[5]), .B(n2610), .Y(n4207) );
  OAI211 U4897 ( .A0(n2611), .A1(n4213), .B0(n4214), .C0(n4215), .Y(N4403) );
  NAND2B U4898 ( .AN(n2745), .B(n4216), .Y(n4215) );
  OAI31 U4899 ( .A0(n2683), .A1(n2602), .A2(n4217), .B0(n4218), .Y(n4216) );
  AOI211 U4900 ( .A0(n2781), .A1(n4219), .B0(n4193), .C0(n4220), .Y(n4214) );
  NOR2 U4901 ( .A(in2_disp[5]), .B(n4188), .Y(n4193) );
  NOR2 U4902 ( .A(n2613), .B(n4204), .Y(n4219) );
  XOR2 U4903 ( .A(in2_disp[5]), .B(n2611), .Y(n4204) );
  AOI22 U4904 ( .A0(n4221), .A1(n2613), .B0(n4198), .B1(in2_disp[5]), .Y(n4213) );
  OAI222 U4905 ( .A0(n4188), .A1(n4222), .B0(n4205), .B1(n4223), .C0(n2746), 
        .C1(n4224), .Y(N4402) );
  NOR2 U4906 ( .A(n2613), .B(in2_disp[5]), .Y(n4222) );
  OAI21 U4907 ( .A0(n4212), .A1(n4205), .B0(n4225), .Y(N4401) );
  AOI211 U4908 ( .A0(n4223), .A1(n4198), .B0(n4226), .C0(n4227), .Y(n4225) );
  NOR2 U4909 ( .A(n4228), .B(n2745), .Y(n4227) );
  INV U4910 ( .A(n4229), .Y(n4226) );
  NAND2B U4911 ( .AN(n2611), .B(n2781), .Y(n4205) );
  OAI211 U4912 ( .A0(n4230), .A1(n2746), .B0(n4231), .C0(n4229), .Y(N4400) );
  NAND2B U4913 ( .AN(n4223), .B(n4221), .Y(n4229) );
  INV U4914 ( .A(n4188), .Y(n4221) );
  NAND2 U4915 ( .A(n2781), .B(in2_disp[7]), .Y(n4188) );
  AOI211 U4916 ( .A0(n4198), .A1(n4232), .B0(n4220), .C0(n4233), .Y(n4231) );
  NOR2B U4917 ( .AN(n4212), .B(n2778), .Y(n4233) );
  NOR2B U4918 ( .AN(in2_disp[5]), .B(n2613), .Y(n4212) );
  NOR3B U4919 ( .AN(n4223), .B(n2777), .C(n2610), .Y(n4220) );
  NOR2B U4920 ( .AN(n2613), .B(in2_disp[5]), .Y(n4223) );
  NOR2B U4921 ( .AN(n2613), .B(n2611), .Y(n4232) );
  NOR2 U4922 ( .A(in2_disp[7]), .B(n2777), .Y(n4198) );
  OAI211 U4923 ( .A0(in2_disp[9]), .A1(n4234), .B0(n4235), .C0(n4236), .Y(
        N4254) );
  AOI2BB2 U4924 ( .B0(n4237), .B1(in2_disp[11]), .A0N(n4238), .A1N(n2745), .Y(
        n4236) );
  AOI211 U4925 ( .A0(in2_disp[10]), .A1(n4239), .B0(n4240), .C0(n4241), .Y(
        n4235) );
  OAI2BB2 U4926 ( .B0(n2780), .B1(n4242), .A0N(in2_disp[8]), .A1N(n4243), .Y(
        n4239) );
  OAI211 U4927 ( .A0(in2_disp[9]), .A1(n4244), .B0(n4245), .C0(n4246), .Y(
        N4253) );
  AOI21 U4928 ( .A0(n4241), .A1(in2_disp[8]), .B0(n4240), .Y(n4246) );
  AOI2BB2 U4929 ( .B0(n4243), .B1(n4247), .A0N(n4248), .A1N(n2746), .Y(n4245)
         );
  NOR2 U4930 ( .A(n4249), .B(n4250), .Y(n4244) );
  NOR2B U4931 ( .AN(n4237), .B(in2_disp[11]), .Y(n4249) );
  OAI211 U4932 ( .A0(n4251), .A1(n2745), .B0(n4252), .C0(n4253), .Y(N4252) );
  OAI2BB1 U4933 ( .A0N(n4254), .A1N(n4255), .B0(n4243), .Y(n4253) );
  NOR2B U4934 ( .AN(n4234), .B(n4256), .Y(n4252) );
  OAI211 U4935 ( .A0(in2_disp[9]), .A1(n4257), .B0(n4258), .C0(n4259), .Y(
        N4251) );
  OAI2BB1 U4936 ( .A0N(n4260), .A1N(n4261), .B0(n4153), .Y(n4259) );
  MX2 U4937 ( .A(n4262), .B(n4263), .S0(in2_disp[10]), .Y(n4258) );
  NOR2 U4938 ( .A(n4256), .B(n4264), .Y(n4263) );
  NOR3 U4939 ( .A(in2_disp[9]), .B(n2779), .C(n4255), .Y(n4256) );
  NOR2 U4940 ( .A(n4241), .B(n4250), .Y(n4262) );
  NOR2B U4941 ( .AN(n4243), .B(n4242), .Y(n4241) );
  NAND2 U4942 ( .A(n4257), .B(n4265), .Y(N4250) );
  AOI211 U4943 ( .A0(n4153), .A1(n4266), .B0(n4267), .C0(n4264), .Y(n4265) );
  NOR2B U4944 ( .AN(n4268), .B(n4242), .Y(n4267) );
  AOI21 U4945 ( .A0(in2_disp[10]), .A1(n4268), .B0(n4240), .Y(n4257) );
  NOR2B U4946 ( .AN(n4237), .B(in2_disp[10]), .Y(n4240) );
  OR2 U4947 ( .A(n4269), .B(n4270), .Y(N4249) );
  OAI222 U4948 ( .A0(n4271), .A1(n4242), .B0(n4272), .B1(n4254), .C0(n2746), 
        .C1(n4273), .Y(n4270) );
  INV U4949 ( .A(n4237), .Y(n4272) );
  INV U4950 ( .A(n4268), .Y(n4271) );
  OAI211 U4951 ( .A0(n4274), .A1(n2745), .B0(n4275), .C0(n4276), .Y(N4248) );
  AOI211 U4952 ( .A0(n2781), .A1(n4254), .B0(n4250), .C0(n4264), .Y(n4276) );
  NOR2B U4953 ( .AN(n4237), .B(n4242), .Y(n4264) );
  NOR2 U4954 ( .A(in2_disp[8]), .B(n2778), .Y(n4237) );
  NOR2B U4955 ( .AN(n4268), .B(n4255), .Y(n4250) );
  INV U4956 ( .A(in2_disp[8]), .Y(n4255) );
  NOR2 U4957 ( .A(in2_disp[10]), .B(n4242), .Y(n4254) );
  INV U4958 ( .A(n4269), .Y(n4275) );
  OAI31 U4959 ( .A0(in2_disp[9]), .A1(n4277), .A2(n4247), .B0(n4234), .Y(n4269) );
  NAND2B U4960 ( .AN(in2_disp[10]), .B(n4268), .Y(n4234) );
  NOR2B U4961 ( .AN(in2_disp[11]), .B(n2777), .Y(n4268) );
  INV U4962 ( .A(n4243), .Y(n4277) );
  NOR2 U4963 ( .A(in2_disp[11]), .B(n2780), .Y(n4243) );
  OAI211 U4964 ( .A0(n2607), .A1(n4278), .B0(n4279), .C0(n4280), .Y(N4102) );
  AOI21 U4965 ( .A0(n4153), .A1(n4281), .B0(n4282), .Y(n4280) );
  MX2 U4966 ( .A(n4283), .B(n4284), .S0(n2609), .Y(n4282) );
  NOR2B U4967 ( .AN(in2_disp[13]), .B(n2779), .Y(n4284) );
  NOR2 U4968 ( .A(n4285), .B(n4286), .Y(n4279) );
  NOR2B U4969 ( .AN(n4287), .B(n4288), .Y(n4286) );
  AOI21 U4970 ( .A0(n2609), .A1(n2607), .B0(in2_disp[13]), .Y(n4288) );
  OAI2BB1 U4971 ( .A0N(n2607), .A1N(n4283), .B0(n4289), .Y(N4101) );
  AOI211 U4972 ( .A0(n4153), .A1(n4290), .B0(n4285), .C0(n4291), .Y(n4289) );
  NOR2B U4973 ( .AN(n4287), .B(n4292), .Y(n4291) );
  NOR2B U4974 ( .AN(n4293), .B(n2608), .Y(n4292) );
  NOR2 U4975 ( .A(n2609), .B(n4294), .Y(n4285) );
  INV U4976 ( .A(n4295), .Y(N4100) );
  AOI211 U4977 ( .A0(n4296), .A1(n2781), .B0(n4297), .C0(n4298), .Y(n4295) );
  OAI22 U4978 ( .A0(n2609), .A1(n4278), .B0(n4299), .B1(n2746), .Y(n4298) );
  NOR2B U4979 ( .AN(n4287), .B(n4300), .Y(n4297) );
  NOR2B U4980 ( .AN(n4301), .B(n2607), .Y(n4300) );
  NOR2 U4981 ( .A(in2_disp[13]), .B(n2606), .Y(n4296) );
  OR4 U4982 ( .A(n4283), .B(n4302), .C(n4303), .D(n4304), .Y(N4099) );
  OAI2BB2 U4983 ( .B0(n2607), .B1(n4305), .A0N(n4153), .A1N(n4306), .Y(n4304)
         );
  OAI31 U4984 ( .A0(n2681), .A1(n2598), .A2(n4307), .B0(n4308), .Y(n4306) );
  AOI22 U4985 ( .A0(n4309), .A1(n2609), .B0(n4287), .B1(in2_disp[13]), .Y(
        n4305) );
  NOR3 U4986 ( .A(n2609), .B(n4293), .C(n2778), .Y(n4302) );
  XOR2 U4987 ( .A(in2_disp[13]), .B(n2607), .Y(n4293) );
  NOR2 U4988 ( .A(in2_disp[13]), .B(n4278), .Y(n4283) );
  OAI222 U4989 ( .A0(n4278), .A1(n4310), .B0(n4294), .B1(n4311), .C0(n2745), 
        .C1(n4312), .Y(N4098) );
  NOR2 U4990 ( .A(n2609), .B(in2_disp[13]), .Y(n4310) );
  OAI21 U4991 ( .A0(n4301), .A1(n4294), .B0(n4313), .Y(N4097) );
  AOI211 U4992 ( .A0(n4311), .A1(n4287), .B0(n4314), .C0(n4315), .Y(n4313) );
  NOR2 U4993 ( .A(n4316), .B(n2746), .Y(n4315) );
  INV U4994 ( .A(n4317), .Y(n4314) );
  NAND2B U4995 ( .AN(n2607), .B(n2781), .Y(n4294) );
  OAI211 U4996 ( .A0(n4318), .A1(n2745), .B0(n4319), .C0(n4317), .Y(N4096) );
  NAND2B U4997 ( .AN(n4311), .B(n4309), .Y(n4317) );
  INV U4998 ( .A(n4278), .Y(n4309) );
  NAND2 U4999 ( .A(n2781), .B(in2_disp[15]), .Y(n4278) );
  AOI211 U5000 ( .A0(n4287), .A1(n4320), .B0(n4303), .C0(n4321), .Y(n4319) );
  NOR2B U5001 ( .AN(n4301), .B(n2777), .Y(n4321) );
  NOR2B U5002 ( .AN(in2_disp[13]), .B(n2609), .Y(n4301) );
  NOR3B U5003 ( .AN(n4311), .B(n2780), .C(n2606), .Y(n4303) );
  NOR2B U5004 ( .AN(n2609), .B(in2_disp[13]), .Y(n4311) );
  NOR2B U5005 ( .AN(n2609), .B(n2607), .Y(n4320) );
  NOR2 U5006 ( .A(in2_disp[15]), .B(n2779), .Y(n4287) );
  NOR2B U5007 ( .AN(n4147), .B(n2778), .Y(N3952) );
  AOI21 U5008 ( .A0(n4322), .A1(n4323), .B0(n4324), .Y(n4147) );
  MX2 U5009 ( .A(n4325), .B(n4326), .S0(n4327), .Y(n4324) );
  NOR2 U5010 ( .A(in2_disp[17]), .B(n2677), .Y(n4326) );
  NOR2B U5011 ( .AN(n4328), .B(n4322), .Y(n4325) );
  NOR2B U5012 ( .AN(n4154), .B(n2777), .Y(N3951) );
  OAI211 U5013 ( .A0(in2_disp[17]), .A1(n4329), .B0(n4330), .C0(n4331), .Y(
        n4154) );
  INV U5014 ( .A(n4332), .Y(n4331) );
  MX2 U5015 ( .A(n4333), .B(n4334), .S0(n2605), .Y(n4330) );
  INV U5016 ( .A(n4328), .Y(n4334) );
  NOR2 U5017 ( .A(n4323), .B(n4171), .Y(n4333) );
  NOR2B U5018 ( .AN(n2677), .B(n4335), .Y(n4323) );
  INV U5019 ( .A(n4336), .Y(n4329) );
  NOR2 U5020 ( .A(n4164), .B(n2780), .Y(N3950) );
  NOR4 U5021 ( .A(n4322), .B(n4327), .C(n4337), .D(n4338), .Y(n4164) );
  NOR2B U5022 ( .AN(n2677), .B(n4339), .Y(n4338) );
  NOR2 U5023 ( .A(n2605), .B(in2_disp[17]), .Y(n4337) );
  NOR2B U5024 ( .AN(n4340), .B(n2779), .Y(N3949) );
  OAI31 U5025 ( .A0(n2677), .A1(n4335), .A2(n4171), .B0(n4172), .Y(n4340) );
  MX2 U5026 ( .A(n4341), .B(n4342), .S0(in2_disp[17]), .Y(n4172) );
  NOR3 U5027 ( .A(n2605), .B(n4332), .C(n4342), .Y(n4341) );
  NOR2 U5028 ( .A(n4336), .B(n4343), .Y(n4342) );
  NOR2B U5029 ( .AN(n2677), .B(in2_disp[18]), .Y(n4343) );
  NOR2 U5030 ( .A(n4177), .B(n2778), .Y(N3948) );
  NOR3B U5031 ( .AN(n4344), .B(n4332), .C(n4339), .Y(n4177) );
  NOR2 U5032 ( .A(in2_disp[18]), .B(n2677), .Y(n4332) );
  AOI22 U5033 ( .A0(in2_disp[18]), .A1(n2605), .B0(in2_disp[17]), .B1(n2676), 
        .Y(n4344) );
  NOR2 U5034 ( .A(n4182), .B(n2777), .Y(N3947) );
  NOR3 U5035 ( .A(n4322), .B(n4339), .C(n4345), .Y(n4182) );
  OAI2BB2 U5036 ( .B0(n2677), .B1(n4346), .A0N(n4327), .A1N(n4335), .Y(n4345)
         );
  NOR2B U5037 ( .AN(in2_disp[18]), .B(n2605), .Y(n4327) );
  NOR2 U5038 ( .A(in2_disp[18]), .B(n4335), .Y(n4346) );
  NOR2B U5039 ( .AN(n2605), .B(n4335), .Y(n4339) );
  NOR2B U5040 ( .AN(n2605), .B(in2_disp[18]), .Y(n4322) );
  NOR2 U5041 ( .A(n4184), .B(n2780), .Y(N3946) );
  NOR2B U5042 ( .AN(n4347), .B(n4348), .Y(n4184) );
  AOI2BB1 U5043 ( .A0N(in2_disp[17]), .A1N(n4171), .B0(n2604), .Y(n4348) );
  MX2 U5044 ( .A(n4335), .B(n4349), .S0(in2_disp[18]), .Y(n4347) );
  NOR2 U5045 ( .A(n4328), .B(n4336), .Y(n4349) );
  NOR2 U5046 ( .A(n2605), .B(n2677), .Y(n4336) );
  NOR2B U5047 ( .AN(n2677), .B(in2_disp[17]), .Y(n4328) );
  NOR2B U5048 ( .AN(n4195), .B(n2779), .Y(N3873) );
  AOI21 U5049 ( .A0(n4350), .A1(n4351), .B0(n4352), .Y(n4195) );
  MX2 U5050 ( .A(n4353), .B(n4354), .S0(n4355), .Y(n4352) );
  NOR2 U5051 ( .A(in2_disp[21]), .B(n2683), .Y(n4354) );
  NOR2B U5052 ( .AN(n4356), .B(n4350), .Y(n4353) );
  NOR2B U5053 ( .AN(n4201), .B(n2778), .Y(N3872) );
  OAI211 U5054 ( .A0(in2_disp[21]), .A1(n4357), .B0(n4358), .C0(n4359), .Y(
        n4201) );
  INV U5055 ( .A(n4360), .Y(n4359) );
  MX2 U5056 ( .A(n4361), .B(n4362), .S0(n2603), .Y(n4358) );
  INV U5057 ( .A(n4356), .Y(n4362) );
  NOR2 U5058 ( .A(n4351), .B(n4217), .Y(n4361) );
  NOR2B U5059 ( .AN(n2683), .B(n4363), .Y(n4351) );
  INV U5060 ( .A(n4364), .Y(n4357) );
  NOR2 U5061 ( .A(n4210), .B(n2777), .Y(N3871) );
  NOR4 U5062 ( .A(n4350), .B(n4355), .C(n4365), .D(n4366), .Y(n4210) );
  NOR2B U5063 ( .AN(n2683), .B(n4367), .Y(n4366) );
  NOR2 U5064 ( .A(n2603), .B(in2_disp[21]), .Y(n4365) );
  NOR2B U5065 ( .AN(n4368), .B(n2780), .Y(N3870) );
  OAI31 U5066 ( .A0(n2683), .A1(n4363), .A2(n4217), .B0(n4218), .Y(n4368) );
  MX2 U5067 ( .A(n4369), .B(n4370), .S0(in2_disp[21]), .Y(n4218) );
  NOR3 U5068 ( .A(n2603), .B(n4360), .C(n4370), .Y(n4369) );
  NOR2 U5069 ( .A(n4364), .B(n4371), .Y(n4370) );
  NOR2B U5070 ( .AN(n2683), .B(in2_disp[22]), .Y(n4371) );
  NOR2 U5071 ( .A(n4224), .B(n2779), .Y(N3869) );
  NOR3B U5072 ( .AN(n4372), .B(n4360), .C(n4367), .Y(n4224) );
  NOR2 U5073 ( .A(in2_disp[22]), .B(n2683), .Y(n4360) );
  AOI22 U5074 ( .A0(in2_disp[22]), .A1(n2603), .B0(in2_disp[21]), .B1(n2682), 
        .Y(n4372) );
  NOR2 U5075 ( .A(n4228), .B(n2778), .Y(N3868) );
  NOR3 U5076 ( .A(n4350), .B(n4367), .C(n4373), .Y(n4228) );
  OAI2BB2 U5077 ( .B0(n2683), .B1(n4374), .A0N(n4355), .A1N(n4363), .Y(n4373)
         );
  NOR2B U5078 ( .AN(in2_disp[22]), .B(n2603), .Y(n4355) );
  NOR2 U5079 ( .A(in2_disp[22]), .B(n4363), .Y(n4374) );
  NOR2B U5080 ( .AN(n2603), .B(n4363), .Y(n4367) );
  NOR2B U5081 ( .AN(n2603), .B(in2_disp[22]), .Y(n4350) );
  NOR2 U5082 ( .A(n4230), .B(n2777), .Y(N3867) );
  NOR2B U5083 ( .AN(n4375), .B(n4376), .Y(n4230) );
  AOI2BB1 U5084 ( .A0N(in2_disp[21]), .A1N(n4217), .B0(n2602), .Y(n4376) );
  MX2 U5085 ( .A(n4363), .B(n4377), .S0(in2_disp[22]), .Y(n4375) );
  NOR2 U5086 ( .A(n4356), .B(n4364), .Y(n4377) );
  NOR2 U5087 ( .A(n2603), .B(n2683), .Y(n4364) );
  NOR2B U5088 ( .AN(n2683), .B(in2_disp[21]), .Y(n4356) );
  NOR2 U5089 ( .A(n4238), .B(n2780), .Y(N3794) );
  NOR4B U5090 ( .AN(n4378), .B(n4379), .C(n4380), .D(n4381), .Y(n4238) );
  MX2 U5091 ( .A(n4382), .B(n4383), .S0(n2601), .Y(n4378) );
  NOR2 U5092 ( .A(in2_disp[25]), .B(n4384), .Y(n4382) );
  NOR2 U5093 ( .A(n4248), .B(n2779), .Y(N3793) );
  AOI211 U5094 ( .A0(n2601), .A1(n4385), .B0(n4386), .C0(n4379), .Y(n4248) );
  AOI211 U5095 ( .A0(in2_disp[24]), .A1(n4387), .B0(n2601), .C0(n4388), .Y(
        n4386) );
  NOR2 U5096 ( .A(in2_disp[25]), .B(n4389), .Y(n4385) );
  NOR2 U5097 ( .A(n4251), .B(n2778), .Y(N3792) );
  AOI211 U5098 ( .A0(n2601), .A1(n4390), .B0(n4391), .C0(n4392), .Y(n4251) );
  NOR2 U5099 ( .A(in2_disp[25]), .B(n4380), .Y(n4392) );
  NOR2 U5100 ( .A(n4393), .B(n2777), .Y(N3791) );
  NOR2B U5101 ( .AN(n4260), .B(n4388), .Y(n4393) );
  NOR2B U5102 ( .AN(n4381), .B(in2_disp[24]), .Y(n4388) );
  MX2 U5103 ( .A(in2_disp[25]), .B(n4394), .S0(n4395), .Y(n4260) );
  NOR2 U5104 ( .A(n4384), .B(n4380), .Y(n4395) );
  NOR2B U5105 ( .AN(in2_disp[26]), .B(n4389), .Y(n4384) );
  NOR2B U5106 ( .AN(n4391), .B(in2_disp[25]), .Y(n4394) );
  NOR2 U5107 ( .A(n2601), .B(n4379), .Y(n4391) );
  NOR2 U5108 ( .A(in2_disp[26]), .B(in2_disp[24]), .Y(n4379) );
  NOR2B U5109 ( .AN(n4266), .B(n2780), .Y(N3790) );
  OAI2BB2 U5110 ( .B0(in2_disp[24]), .B1(n4387), .A0N(n2601), .A1N(n4383), .Y(
        n4266) );
  NOR2 U5111 ( .A(n4273), .B(n2779), .Y(N3789) );
  AOI211 U5112 ( .A0(n4387), .A1(n2600), .B0(n4396), .C0(n4397), .Y(n4273) );
  AOI21 U5113 ( .A0(in2_disp[25]), .A1(n4390), .B0(in2_disp[24]), .Y(n4396) );
  NOR2 U5114 ( .A(n4274), .B(n2778), .Y(N3788) );
  NOR2B U5115 ( .AN(n4398), .B(n4397), .Y(n4274) );
  NOR2B U5116 ( .AN(n2601), .B(n4387), .Y(n4397) );
  NOR2 U5117 ( .A(in2_disp[25]), .B(n4390), .Y(n4387) );
  OAI211 U5118 ( .A0(n4389), .A1(n4399), .B0(n4383), .C0(n4261), .Y(n4398) );
  NAND2 U5119 ( .A(in2_disp[26]), .B(n4380), .Y(n4261) );
  NOR2B U5120 ( .AN(n2601), .B(in2_disp[24]), .Y(n4380) );
  OR2 U5121 ( .A(in2_disp[26]), .B(in2_disp[25]), .Y(n4383) );
  INV U5122 ( .A(n4381), .Y(n4399) );
  NOR2B U5123 ( .AN(in2_disp[25]), .B(n4390), .Y(n4381) );
  INV U5124 ( .A(in2_disp[24]), .Y(n4389) );
  NOR2B U5125 ( .AN(n4281), .B(n2777), .Y(N3715) );
  AOI21 U5126 ( .A0(n4400), .A1(n4401), .B0(n4402), .Y(n4281) );
  MX2 U5127 ( .A(n4403), .B(n4404), .S0(n4405), .Y(n4402) );
  NOR2 U5128 ( .A(in2_disp[29]), .B(n2681), .Y(n4404) );
  NOR2B U5129 ( .AN(n4406), .B(n4400), .Y(n4403) );
  NOR2B U5130 ( .AN(n4290), .B(n2780), .Y(N3714) );
  OAI211 U5131 ( .A0(in2_disp[29]), .A1(n4407), .B0(n4408), .C0(n4409), .Y(
        n4290) );
  INV U5132 ( .A(n4410), .Y(n4409) );
  MX2 U5133 ( .A(n4411), .B(n4412), .S0(n2599), .Y(n4408) );
  INV U5134 ( .A(n4406), .Y(n4412) );
  NOR2 U5135 ( .A(n4401), .B(n4307), .Y(n4411) );
  NOR2B U5136 ( .AN(n2681), .B(n4413), .Y(n4401) );
  INV U5137 ( .A(n4414), .Y(n4407) );
  NOR2 U5138 ( .A(n4299), .B(n2779), .Y(N3713) );
  NOR4 U5139 ( .A(n4400), .B(n4405), .C(n4415), .D(n4416), .Y(n4299) );
  NOR2B U5140 ( .AN(n2681), .B(n4417), .Y(n4416) );
  NOR2 U5141 ( .A(n2599), .B(in2_disp[29]), .Y(n4415) );
  NOR2B U5142 ( .AN(n4418), .B(n2778), .Y(N3712) );
  OAI31 U5143 ( .A0(n2681), .A1(n4413), .A2(n4307), .B0(n4308), .Y(n4418) );
  MX2 U5144 ( .A(n4419), .B(n4420), .S0(in2_disp[29]), .Y(n4308) );
  NOR3 U5145 ( .A(n2599), .B(n4410), .C(n4420), .Y(n4419) );
  NOR2 U5146 ( .A(n4414), .B(n4421), .Y(n4420) );
  NOR2B U5147 ( .AN(n2681), .B(in2_disp[30]), .Y(n4421) );
  NOR2 U5148 ( .A(n4312), .B(n2777), .Y(N3711) );
  NOR3B U5149 ( .AN(n4422), .B(n4410), .C(n4417), .Y(n4312) );
  NOR2 U5150 ( .A(in2_disp[30]), .B(n2681), .Y(n4410) );
  AOI22 U5151 ( .A0(in2_disp[30]), .A1(n2599), .B0(in2_disp[29]), .B1(n2680), 
        .Y(n4422) );
  NOR2 U5152 ( .A(n4316), .B(n2780), .Y(N3710) );
  NOR3 U5153 ( .A(n4400), .B(n4417), .C(n4423), .Y(n4316) );
  OAI2BB2 U5154 ( .B0(n2681), .B1(n4424), .A0N(n4405), .A1N(n4413), .Y(n4423)
         );
  NOR2B U5155 ( .AN(in2_disp[30]), .B(n2599), .Y(n4405) );
  NOR2 U5156 ( .A(in2_disp[30]), .B(n4413), .Y(n4424) );
  NOR2B U5157 ( .AN(n2599), .B(n4413), .Y(n4417) );
  NOR2B U5158 ( .AN(n2599), .B(in2_disp[30]), .Y(n4400) );
  NOR2 U5159 ( .A(n4318), .B(n2779), .Y(N3709) );
  NOR2B U5160 ( .AN(n4425), .B(n4426), .Y(n4318) );
  AOI2BB1 U5161 ( .A0N(in2_disp[29]), .A1N(n4307), .B0(n2598), .Y(n4426) );
  MX2 U5162 ( .A(n4413), .B(n4427), .S0(in2_disp[30]), .Y(n4425) );
  NOR2 U5163 ( .A(n4406), .B(n4414), .Y(n4427) );
  NOR2 U5164 ( .A(n2599), .B(n2681), .Y(n4414) );
  NOR2B U5165 ( .AN(n2681), .B(in2_disp[29]), .Y(n4406) );
  OAI211 U5166 ( .A0(n2635), .A1(n4428), .B0(n4429), .C0(n4430), .Y(N3634) );
  AOI21 U5167 ( .A0(n4153), .A1(n4431), .B0(n4432), .Y(n4430) );
  MX2 U5168 ( .A(n4433), .B(n4434), .S0(n2637), .Y(n4432) );
  NOR2B U5169 ( .AN(in1_disp[1]), .B(n2778), .Y(n4434) );
  NOR2 U5170 ( .A(n4435), .B(n4436), .Y(n4429) );
  NOR2B U5171 ( .AN(n4437), .B(n4438), .Y(n4436) );
  AOI21 U5172 ( .A0(n2637), .A1(n2635), .B0(in1_disp[1]), .Y(n4438) );
  OAI2BB1 U5173 ( .A0N(n2635), .A1N(n4433), .B0(n4439), .Y(N3633) );
  AOI211 U5174 ( .A0(n4153), .A1(n4440), .B0(n4435), .C0(n4441), .Y(n4439) );
  NOR2B U5175 ( .AN(n4437), .B(n4442), .Y(n4441) );
  NOR2B U5176 ( .AN(n4443), .B(n2636), .Y(n4442) );
  NOR2 U5177 ( .A(n2637), .B(n4444), .Y(n4435) );
  INV U5178 ( .A(n4445), .Y(N3632) );
  AOI211 U5179 ( .A0(n4446), .A1(n2781), .B0(n4447), .C0(n4448), .Y(n4445) );
  OAI22 U5180 ( .A0(n2637), .A1(n4428), .B0(n4449), .B1(n2746), .Y(n4448) );
  NOR2B U5181 ( .AN(n4437), .B(n4450), .Y(n4447) );
  NOR2B U5182 ( .AN(n4451), .B(n2635), .Y(n4450) );
  NOR2 U5183 ( .A(in1_disp[1]), .B(n2634), .Y(n4446) );
  OR4 U5184 ( .A(n4433), .B(n4452), .C(n4453), .D(n4454), .Y(N3631) );
  OAI2BB2 U5185 ( .B0(n2635), .B1(n4455), .A0N(n4153), .A1N(n4456), .Y(n4454)
         );
  OAI31 U5186 ( .A0(n2675), .A1(n2624), .A2(n4457), .B0(n4458), .Y(n4456) );
  AOI22 U5187 ( .A0(n4459), .A1(n2637), .B0(n4437), .B1(in1_disp[1]), .Y(n4455) );
  NOR3 U5188 ( .A(n2637), .B(n4443), .C(n2777), .Y(n4452) );
  XOR2 U5189 ( .A(in1_disp[1]), .B(n2635), .Y(n4443) );
  NOR2 U5190 ( .A(in1_disp[1]), .B(n4428), .Y(n4433) );
  OAI222 U5191 ( .A0(n4428), .A1(n4460), .B0(n4444), .B1(n4461), .C0(n2745), 
        .C1(n4462), .Y(N3630) );
  NOR2 U5192 ( .A(n2637), .B(in1_disp[1]), .Y(n4460) );
  OAI21 U5193 ( .A0(n4451), .A1(n4444), .B0(n4463), .Y(N3629) );
  AOI211 U5194 ( .A0(n4461), .A1(n4437), .B0(n4464), .C0(n4465), .Y(n4463) );
  NOR2 U5195 ( .A(n4466), .B(n2746), .Y(n4465) );
  INV U5196 ( .A(n4467), .Y(n4464) );
  NAND2B U5197 ( .AN(n2635), .B(n2781), .Y(n4444) );
  OAI211 U5198 ( .A0(n4468), .A1(n2745), .B0(n4469), .C0(n4467), .Y(N3628) );
  NAND2B U5199 ( .AN(n4461), .B(n4459), .Y(n4467) );
  INV U5200 ( .A(n4428), .Y(n4459) );
  NAND2 U5201 ( .A(n2781), .B(in1_disp[3]), .Y(n4428) );
  AOI211 U5202 ( .A0(n4437), .A1(n4470), .B0(n4453), .C0(n4471), .Y(n4469) );
  NOR2B U5203 ( .AN(n4451), .B(n2780), .Y(n4471) );
  NOR2B U5204 ( .AN(in1_disp[1]), .B(n2637), .Y(n4451) );
  NOR3B U5205 ( .AN(n4461), .B(n2779), .C(n2634), .Y(n4453) );
  NOR2B U5206 ( .AN(n2637), .B(in1_disp[1]), .Y(n4461) );
  NOR2B U5207 ( .AN(n2637), .B(n2635), .Y(n4470) );
  NOR2 U5208 ( .A(in1_disp[3]), .B(n2778), .Y(n4437) );
  OAI211 U5209 ( .A0(n2631), .A1(n4472), .B0(n4473), .C0(n4474), .Y(N3482) );
  AOI21 U5210 ( .A0(n4153), .A1(n4475), .B0(n4476), .Y(n4474) );
  MX2 U5211 ( .A(n4477), .B(n4478), .S0(n2633), .Y(n4476) );
  NOR2B U5212 ( .AN(in1_disp[5]), .B(n2777), .Y(n4478) );
  NOR2 U5213 ( .A(n4479), .B(n4480), .Y(n4473) );
  NOR2B U5214 ( .AN(n4481), .B(n4482), .Y(n4480) );
  AOI21 U5215 ( .A0(n2633), .A1(n2631), .B0(in1_disp[5]), .Y(n4482) );
  OAI2BB1 U5216 ( .A0N(n2631), .A1N(n4477), .B0(n4483), .Y(N3481) );
  AOI211 U5217 ( .A0(n4153), .A1(n4484), .B0(n4479), .C0(n4485), .Y(n4483) );
  NOR2B U5218 ( .AN(n4481), .B(n4486), .Y(n4485) );
  NOR2B U5219 ( .AN(n4487), .B(n2632), .Y(n4486) );
  NOR2 U5220 ( .A(n2633), .B(n4488), .Y(n4479) );
  INV U5221 ( .A(n4489), .Y(N3480) );
  AOI211 U5222 ( .A0(n4490), .A1(n2781), .B0(n4491), .C0(n4492), .Y(n4489) );
  OAI22 U5223 ( .A0(n2633), .A1(n4472), .B0(n4493), .B1(n2746), .Y(n4492) );
  NOR2B U5224 ( .AN(n4481), .B(n4494), .Y(n4491) );
  NOR2B U5225 ( .AN(n4495), .B(n2631), .Y(n4494) );
  NOR2 U5226 ( .A(in1_disp[5]), .B(n2630), .Y(n4490) );
  OR4 U5227 ( .A(n4477), .B(n4496), .C(n4497), .D(n4498), .Y(N3479) );
  OAI2BB2 U5228 ( .B0(n2631), .B1(n4499), .A0N(n4153), .A1N(n4500), .Y(n4498)
         );
  OAI31 U5229 ( .A0(n2673), .A1(n2622), .A2(n4501), .B0(n4502), .Y(n4500) );
  AOI22 U5230 ( .A0(n4503), .A1(n2633), .B0(n4481), .B1(in1_disp[5]), .Y(n4499) );
  NOR3 U5231 ( .A(n2633), .B(n4487), .C(n2780), .Y(n4496) );
  XOR2 U5232 ( .A(in1_disp[5]), .B(n2631), .Y(n4487) );
  NOR2 U5233 ( .A(in1_disp[5]), .B(n4472), .Y(n4477) );
  OAI222 U5234 ( .A0(n4472), .A1(n4504), .B0(n4488), .B1(n4505), .C0(n2745), 
        .C1(n4506), .Y(N3478) );
  NOR2 U5235 ( .A(n2633), .B(in1_disp[5]), .Y(n4504) );
  OAI21 U5236 ( .A0(n4495), .A1(n4488), .B0(n4507), .Y(N3477) );
  AOI211 U5237 ( .A0(n4505), .A1(n4481), .B0(n4508), .C0(n4509), .Y(n4507) );
  NOR2 U5238 ( .A(n4510), .B(n2746), .Y(n4509) );
  INV U5239 ( .A(n4511), .Y(n4508) );
  NAND2B U5240 ( .AN(n2631), .B(n2781), .Y(n4488) );
  OAI211 U5241 ( .A0(n4512), .A1(n2745), .B0(n4513), .C0(n4511), .Y(N3476) );
  NAND2B U5242 ( .AN(n4505), .B(n4503), .Y(n4511) );
  INV U5243 ( .A(n4472), .Y(n4503) );
  NAND2 U5244 ( .A(n2781), .B(in1_disp[7]), .Y(n4472) );
  AOI211 U5245 ( .A0(n4481), .A1(n4514), .B0(n4497), .C0(n4515), .Y(n4513) );
  NOR2B U5246 ( .AN(n4495), .B(n2779), .Y(n4515) );
  NOR2B U5247 ( .AN(in1_disp[5]), .B(n2633), .Y(n4495) );
  NOR3B U5248 ( .AN(n4505), .B(n2778), .C(n2630), .Y(n4497) );
  NOR2B U5249 ( .AN(n2633), .B(in1_disp[5]), .Y(n4505) );
  NOR2B U5250 ( .AN(n2633), .B(n2631), .Y(n4514) );
  NOR2 U5251 ( .A(in1_disp[7]), .B(n2777), .Y(n4481) );
  OAI211 U5252 ( .A0(in1_disp[9]), .A1(n4516), .B0(n4517), .C0(n4518), .Y(
        N3330) );
  AOI2BB2 U5253 ( .B0(n4519), .B1(in1_disp[11]), .A0N(n4520), .A1N(n2746), .Y(
        n4518) );
  AOI211 U5254 ( .A0(in1_disp[10]), .A1(n4521), .B0(n4522), .C0(n4523), .Y(
        n4517) );
  OAI2BB2 U5255 ( .B0(n2780), .B1(n4524), .A0N(in1_disp[8]), .A1N(n4525), .Y(
        n4521) );
  OAI211 U5256 ( .A0(in1_disp[9]), .A1(n4526), .B0(n4527), .C0(n4528), .Y(
        N3329) );
  AOI21 U5257 ( .A0(n4523), .A1(in1_disp[8]), .B0(n4522), .Y(n4528) );
  AOI2BB2 U5258 ( .B0(n4525), .B1(n4529), .A0N(n4530), .A1N(n2745), .Y(n4527)
         );
  NOR2 U5259 ( .A(n4531), .B(n4532), .Y(n4526) );
  NOR2B U5260 ( .AN(n4519), .B(in1_disp[11]), .Y(n4531) );
  OAI211 U5261 ( .A0(n4533), .A1(n2746), .B0(n4534), .C0(n4535), .Y(N3328) );
  OAI2BB1 U5262 ( .A0N(n4536), .A1N(n4537), .B0(n4525), .Y(n4535) );
  NOR2B U5263 ( .AN(n4516), .B(n4538), .Y(n4534) );
  OAI211 U5264 ( .A0(in1_disp[9]), .A1(n4539), .B0(n4540), .C0(n4541), .Y(
        N3327) );
  OAI2BB1 U5265 ( .A0N(n4542), .A1N(n4543), .B0(n4153), .Y(n4541) );
  MX2 U5266 ( .A(n4544), .B(n4545), .S0(in1_disp[10]), .Y(n4540) );
  NOR2 U5267 ( .A(n4538), .B(n4546), .Y(n4545) );
  NOR3 U5268 ( .A(in1_disp[9]), .B(n2779), .C(n4537), .Y(n4538) );
  NOR2 U5269 ( .A(n4523), .B(n4532), .Y(n4544) );
  NOR2B U5270 ( .AN(n4525), .B(n4524), .Y(n4523) );
  NAND2 U5271 ( .A(n4539), .B(n4547), .Y(N3326) );
  AOI211 U5272 ( .A0(n4153), .A1(n4548), .B0(n4549), .C0(n4546), .Y(n4547) );
  NOR2B U5273 ( .AN(n4550), .B(n4524), .Y(n4549) );
  AOI21 U5274 ( .A0(in1_disp[10]), .A1(n4550), .B0(n4522), .Y(n4539) );
  NOR2B U5275 ( .AN(n4519), .B(in1_disp[10]), .Y(n4522) );
  OR2 U5276 ( .A(n4551), .B(n4552), .Y(N3325) );
  OAI222 U5277 ( .A0(n4553), .A1(n4524), .B0(n4554), .B1(n4536), .C0(n2745), 
        .C1(n4555), .Y(n4552) );
  INV U5278 ( .A(n4519), .Y(n4554) );
  INV U5279 ( .A(n4550), .Y(n4553) );
  OAI211 U5280 ( .A0(n4556), .A1(n2746), .B0(n4557), .C0(n4558), .Y(N3324) );
  AOI211 U5281 ( .A0(n2781), .A1(n4536), .B0(n4532), .C0(n4546), .Y(n4558) );
  NOR2B U5282 ( .AN(n4519), .B(n4524), .Y(n4546) );
  NOR2 U5283 ( .A(in1_disp[8]), .B(n2778), .Y(n4519) );
  NOR2B U5284 ( .AN(n4550), .B(n4537), .Y(n4532) );
  INV U5285 ( .A(in1_disp[8]), .Y(n4537) );
  NOR2 U5286 ( .A(in1_disp[10]), .B(n4524), .Y(n4536) );
  INV U5287 ( .A(n4551), .Y(n4557) );
  OAI31 U5288 ( .A0(in1_disp[9]), .A1(n4559), .A2(n4529), .B0(n4516), .Y(n4551) );
  NAND2B U5289 ( .AN(in1_disp[10]), .B(n4550), .Y(n4516) );
  NOR2B U5290 ( .AN(in1_disp[11]), .B(n2777), .Y(n4550) );
  INV U5291 ( .A(n4525), .Y(n4559) );
  NOR2 U5292 ( .A(in1_disp[11]), .B(n2780), .Y(n4525) );
  OAI211 U5293 ( .A0(n2627), .A1(n4560), .B0(n4561), .C0(n4562), .Y(N3178) );
  AOI21 U5294 ( .A0(n4153), .A1(n4563), .B0(n4564), .Y(n4562) );
  MX2 U5295 ( .A(n4565), .B(n4566), .S0(n2629), .Y(n4564) );
  NOR2B U5296 ( .AN(in1_disp[13]), .B(n2779), .Y(n4566) );
  NOR2 U5297 ( .A(n4567), .B(n4568), .Y(n4561) );
  NOR2B U5298 ( .AN(n4569), .B(n4570), .Y(n4568) );
  AOI21 U5299 ( .A0(n2629), .A1(n2627), .B0(in1_disp[13]), .Y(n4570) );
  OAI2BB1 U5300 ( .A0N(n2627), .A1N(n4565), .B0(n4571), .Y(N3177) );
  AOI211 U5301 ( .A0(n4153), .A1(n4572), .B0(n4567), .C0(n4573), .Y(n4571) );
  NOR2B U5302 ( .AN(n4569), .B(n4574), .Y(n4573) );
  NOR2B U5303 ( .AN(n4575), .B(n2628), .Y(n4574) );
  NOR2 U5304 ( .A(n2629), .B(n4576), .Y(n4567) );
  INV U5305 ( .A(n4577), .Y(N3176) );
  AOI211 U5306 ( .A0(n4578), .A1(n2781), .B0(n4579), .C0(n4580), .Y(n4577) );
  OAI22 U5307 ( .A0(n2629), .A1(n4560), .B0(n4581), .B1(n2745), .Y(n4580) );
  NOR2B U5308 ( .AN(n4569), .B(n4582), .Y(n4579) );
  NOR2B U5309 ( .AN(n4583), .B(n2627), .Y(n4582) );
  NOR2 U5310 ( .A(in1_disp[13]), .B(n2626), .Y(n4578) );
  OR4 U5311 ( .A(n4565), .B(n4584), .C(n4585), .D(n4586), .Y(N3175) );
  OAI2BB2 U5312 ( .B0(n2627), .B1(n4587), .A0N(n4153), .A1N(n4588), .Y(n4586)
         );
  OAI31 U5313 ( .A0(n2679), .A1(n2618), .A2(n4589), .B0(n4590), .Y(n4588) );
  INV U5314 ( .A(n2745), .Y(n4153) );
  AOI22 U5315 ( .A0(n4591), .A1(n2629), .B0(n4569), .B1(in1_disp[13]), .Y(
        n4587) );
  NOR3 U5316 ( .A(n2629), .B(n4575), .C(n2778), .Y(n4584) );
  XOR2 U5317 ( .A(in1_disp[13]), .B(n2627), .Y(n4575) );
  NOR2 U5318 ( .A(in1_disp[13]), .B(n4560), .Y(n4565) );
  OAI222 U5319 ( .A0(n4560), .A1(n4592), .B0(n4576), .B1(n4593), .C0(n2746), 
        .C1(n4594), .Y(N3174) );
  NOR2 U5320 ( .A(n2629), .B(in1_disp[13]), .Y(n4592) );
  OAI21 U5321 ( .A0(n4583), .A1(n4576), .B0(n4595), .Y(N3173) );
  AOI211 U5322 ( .A0(n4593), .A1(n4569), .B0(n4596), .C0(n4597), .Y(n4595) );
  NOR2 U5323 ( .A(n4598), .B(n2745), .Y(n4597) );
  INV U5324 ( .A(n4599), .Y(n4596) );
  NAND2B U5325 ( .AN(n2627), .B(n2781), .Y(n4576) );
  OAI211 U5326 ( .A0(n4600), .A1(n2746), .B0(n4601), .C0(n4599), .Y(N3172) );
  NAND2B U5327 ( .AN(n4593), .B(n4591), .Y(n4599) );
  INV U5328 ( .A(n4560), .Y(n4591) );
  NAND2 U5329 ( .A(n2781), .B(in1_disp[15]), .Y(n4560) );
  AOI211 U5330 ( .A0(n4569), .A1(n4602), .B0(n4585), .C0(n4603), .Y(n4601) );
  NOR2B U5331 ( .AN(n4583), .B(n2777), .Y(n4603) );
  NOR2B U5332 ( .AN(in1_disp[13]), .B(n2629), .Y(n4583) );
  NOR3B U5333 ( .AN(n4593), .B(n2780), .C(n2626), .Y(n4585) );
  NOR2B U5334 ( .AN(n2629), .B(in1_disp[13]), .Y(n4593) );
  NOR2B U5335 ( .AN(n2629), .B(n2627), .Y(n4602) );
  NOR2 U5336 ( .A(in1_disp[15]), .B(n2779), .Y(n4569) );
  NOR2B U5337 ( .AN(n4431), .B(n2778), .Y(N3028) );
  AOI21 U5338 ( .A0(n4604), .A1(n4605), .B0(n4606), .Y(n4431) );
  MX2 U5339 ( .A(n4607), .B(n4608), .S0(n4609), .Y(n4606) );
  NOR2 U5340 ( .A(in1_disp[17]), .B(n2675), .Y(n4608) );
  NOR2B U5341 ( .AN(n4610), .B(n4604), .Y(n4607) );
  NOR2B U5342 ( .AN(n4440), .B(n2777), .Y(N3027) );
  OAI211 U5343 ( .A0(in1_disp[17]), .A1(n4611), .B0(n4612), .C0(n4613), .Y(
        n4440) );
  INV U5344 ( .A(n4614), .Y(n4613) );
  MX2 U5345 ( .A(n4615), .B(n4616), .S0(n2625), .Y(n4612) );
  INV U5346 ( .A(n4610), .Y(n4616) );
  NOR2 U5347 ( .A(n4605), .B(n4457), .Y(n4615) );
  NOR2B U5348 ( .AN(n2675), .B(n4617), .Y(n4605) );
  INV U5349 ( .A(n4618), .Y(n4611) );
  NOR2 U5350 ( .A(n4449), .B(n2780), .Y(N3026) );
  NOR4 U5351 ( .A(n4604), .B(n4609), .C(n4619), .D(n4620), .Y(n4449) );
  NOR2B U5352 ( .AN(n2675), .B(n4621), .Y(n4620) );
  NOR2 U5353 ( .A(n2625), .B(in1_disp[17]), .Y(n4619) );
  NOR2B U5354 ( .AN(n4622), .B(n2779), .Y(N3025) );
  OAI31 U5355 ( .A0(n2675), .A1(n4617), .A2(n4457), .B0(n4458), .Y(n4622) );
  MX2 U5356 ( .A(n4623), .B(n4624), .S0(in1_disp[17]), .Y(n4458) );
  NOR3 U5357 ( .A(n2625), .B(n4614), .C(n4624), .Y(n4623) );
  NOR2 U5358 ( .A(n4618), .B(n4625), .Y(n4624) );
  NOR2B U5359 ( .AN(n2675), .B(in1_disp[18]), .Y(n4625) );
  NOR2 U5360 ( .A(n4462), .B(n2778), .Y(N3024) );
  NOR3B U5361 ( .AN(n4626), .B(n4614), .C(n4621), .Y(n4462) );
  NOR2 U5362 ( .A(in1_disp[18]), .B(n2675), .Y(n4614) );
  AOI22 U5363 ( .A0(in1_disp[18]), .A1(n2625), .B0(in1_disp[17]), .B1(n2674), 
        .Y(n4626) );
  NOR2 U5364 ( .A(n4466), .B(n2777), .Y(N3023) );
  NOR3 U5365 ( .A(n4604), .B(n4621), .C(n4627), .Y(n4466) );
  OAI2BB2 U5366 ( .B0(n2675), .B1(n4628), .A0N(n4609), .A1N(n4617), .Y(n4627)
         );
  NOR2B U5367 ( .AN(in1_disp[18]), .B(n2625), .Y(n4609) );
  NOR2 U5368 ( .A(in1_disp[18]), .B(n4617), .Y(n4628) );
  NOR2B U5369 ( .AN(n2625), .B(n4617), .Y(n4621) );
  NOR2B U5370 ( .AN(n2625), .B(in1_disp[18]), .Y(n4604) );
  NOR2 U5371 ( .A(n4468), .B(n2780), .Y(N3022) );
  NOR2B U5372 ( .AN(n4629), .B(n4630), .Y(n4468) );
  AOI2BB1 U5373 ( .A0N(in1_disp[17]), .A1N(n4457), .B0(n2624), .Y(n4630) );
  MX2 U5374 ( .A(n4617), .B(n4631), .S0(in1_disp[18]), .Y(n4629) );
  NOR2 U5375 ( .A(n4610), .B(n4618), .Y(n4631) );
  NOR2 U5376 ( .A(n2625), .B(n2675), .Y(n4618) );
  NOR2B U5377 ( .AN(n2675), .B(in1_disp[17]), .Y(n4610) );
  NOR2B U5378 ( .AN(n4475), .B(n2779), .Y(N2949) );
  AOI21 U5379 ( .A0(n4632), .A1(n4633), .B0(n4634), .Y(n4475) );
  MX2 U5380 ( .A(n4635), .B(n4636), .S0(n4637), .Y(n4634) );
  NOR2 U5381 ( .A(in1_disp[21]), .B(n2673), .Y(n4636) );
  NOR2B U5382 ( .AN(n4638), .B(n4632), .Y(n4635) );
  NOR2B U5383 ( .AN(n4484), .B(n2778), .Y(N2948) );
  OAI211 U5384 ( .A0(in1_disp[21]), .A1(n4639), .B0(n4640), .C0(n4641), .Y(
        n4484) );
  INV U5385 ( .A(n4642), .Y(n4641) );
  MX2 U5386 ( .A(n4643), .B(n4644), .S0(n2623), .Y(n4640) );
  INV U5387 ( .A(n4638), .Y(n4644) );
  NOR2 U5388 ( .A(n4633), .B(n4501), .Y(n4643) );
  NOR2B U5389 ( .AN(n2673), .B(n4645), .Y(n4633) );
  INV U5390 ( .A(n4646), .Y(n4639) );
  NOR2 U5391 ( .A(n4493), .B(n2777), .Y(N2947) );
  NOR4 U5392 ( .A(n4632), .B(n4637), .C(n4647), .D(n4648), .Y(n4493) );
  NOR2B U5393 ( .AN(n2673), .B(n4649), .Y(n4648) );
  NOR2 U5394 ( .A(n2623), .B(in1_disp[21]), .Y(n4647) );
  NOR2B U5395 ( .AN(n4650), .B(n2780), .Y(N2946) );
  OAI31 U5396 ( .A0(n2673), .A1(n4645), .A2(n4501), .B0(n4502), .Y(n4650) );
  MX2 U5397 ( .A(n4651), .B(n4652), .S0(in1_disp[21]), .Y(n4502) );
  NOR3 U5398 ( .A(n2623), .B(n4642), .C(n4652), .Y(n4651) );
  NOR2 U5399 ( .A(n4646), .B(n4653), .Y(n4652) );
  NOR2B U5400 ( .AN(n2673), .B(in1_disp[22]), .Y(n4653) );
  NOR2 U5401 ( .A(n4506), .B(n2779), .Y(N2945) );
  NOR3B U5402 ( .AN(n4654), .B(n4642), .C(n4649), .Y(n4506) );
  NOR2 U5403 ( .A(in1_disp[22]), .B(n2673), .Y(n4642) );
  AOI22 U5404 ( .A0(in1_disp[22]), .A1(n2623), .B0(in1_disp[21]), .B1(n2672), 
        .Y(n4654) );
  NOR2 U5405 ( .A(n4510), .B(n2778), .Y(N2944) );
  NOR3 U5406 ( .A(n4632), .B(n4649), .C(n4655), .Y(n4510) );
  OAI2BB2 U5407 ( .B0(n2673), .B1(n4656), .A0N(n4637), .A1N(n4645), .Y(n4655)
         );
  NOR2B U5408 ( .AN(in1_disp[22]), .B(n2623), .Y(n4637) );
  NOR2 U5409 ( .A(in1_disp[22]), .B(n4645), .Y(n4656) );
  NOR2B U5410 ( .AN(n2623), .B(n4645), .Y(n4649) );
  NOR2B U5411 ( .AN(n2623), .B(in1_disp[22]), .Y(n4632) );
  NOR2 U5412 ( .A(n4512), .B(n2777), .Y(N2943) );
  NOR2B U5413 ( .AN(n4657), .B(n4658), .Y(n4512) );
  AOI2BB1 U5414 ( .A0N(in1_disp[21]), .A1N(n4501), .B0(n2622), .Y(n4658) );
  MX2 U5415 ( .A(n4645), .B(n4659), .S0(in1_disp[22]), .Y(n4657) );
  NOR2 U5416 ( .A(n4638), .B(n4646), .Y(n4659) );
  NOR2 U5417 ( .A(n2623), .B(n2673), .Y(n4646) );
  NOR2B U5418 ( .AN(n2673), .B(in1_disp[21]), .Y(n4638) );
  NOR2 U5419 ( .A(n4520), .B(n2780), .Y(N2870) );
  NOR4B U5420 ( .AN(n4660), .B(n4661), .C(n4662), .D(n4663), .Y(n4520) );
  MX2 U5421 ( .A(n4664), .B(n4665), .S0(n2621), .Y(n4660) );
  NOR2 U5422 ( .A(in1_disp[25]), .B(n4666), .Y(n4664) );
  NOR2 U5423 ( .A(n4530), .B(n2779), .Y(N2869) );
  AOI211 U5424 ( .A0(n2621), .A1(n4667), .B0(n4668), .C0(n4661), .Y(n4530) );
  AOI211 U5425 ( .A0(in1_disp[24]), .A1(n4669), .B0(n2621), .C0(n4670), .Y(
        n4668) );
  NOR2 U5426 ( .A(in1_disp[25]), .B(n4671), .Y(n4667) );
  NOR2 U5427 ( .A(n4533), .B(n2778), .Y(N2868) );
  AOI211 U5428 ( .A0(n2621), .A1(n4672), .B0(n4673), .C0(n4674), .Y(n4533) );
  NOR2 U5429 ( .A(in1_disp[25]), .B(n4662), .Y(n4674) );
  NOR2 U5430 ( .A(n4675), .B(n2777), .Y(N2867) );
  NOR2B U5431 ( .AN(n4542), .B(n4670), .Y(n4675) );
  NOR2B U5432 ( .AN(n4663), .B(in1_disp[24]), .Y(n4670) );
  MX2 U5433 ( .A(in1_disp[25]), .B(n4676), .S0(n4677), .Y(n4542) );
  NOR2 U5434 ( .A(n4666), .B(n4662), .Y(n4677) );
  NOR2B U5435 ( .AN(in1_disp[26]), .B(n4671), .Y(n4666) );
  NOR2B U5436 ( .AN(n4673), .B(in1_disp[25]), .Y(n4676) );
  NOR2 U5437 ( .A(n2621), .B(n4661), .Y(n4673) );
  NOR2 U5438 ( .A(in1_disp[26]), .B(in1_disp[24]), .Y(n4661) );
  NOR2B U5439 ( .AN(n4548), .B(n2780), .Y(N2866) );
  OAI2BB2 U5440 ( .B0(in1_disp[24]), .B1(n4669), .A0N(n2621), .A1N(n4665), .Y(
        n4548) );
  NOR2 U5441 ( .A(n4555), .B(n2779), .Y(N2865) );
  AOI211 U5442 ( .A0(n4669), .A1(n2620), .B0(n4678), .C0(n4679), .Y(n4555) );
  AOI21 U5443 ( .A0(in1_disp[25]), .A1(n4672), .B0(in1_disp[24]), .Y(n4678) );
  NOR2 U5444 ( .A(n4556), .B(n2778), .Y(N2864) );
  NOR2B U5445 ( .AN(n4680), .B(n4679), .Y(n4556) );
  NOR2B U5446 ( .AN(n2621), .B(n4669), .Y(n4679) );
  NOR2 U5447 ( .A(in1_disp[25]), .B(n4672), .Y(n4669) );
  OAI211 U5448 ( .A0(n4671), .A1(n4681), .B0(n4665), .C0(n4543), .Y(n4680) );
  NAND2 U5449 ( .A(in1_disp[26]), .B(n4662), .Y(n4543) );
  NOR2B U5450 ( .AN(n2621), .B(in1_disp[24]), .Y(n4662) );
  OR2 U5451 ( .A(in1_disp[26]), .B(in1_disp[25]), .Y(n4665) );
  INV U5452 ( .A(n4663), .Y(n4681) );
  NOR2B U5453 ( .AN(in1_disp[25]), .B(n4672), .Y(n4663) );
  INV U5454 ( .A(in1_disp[24]), .Y(n4671) );
  NOR2B U5455 ( .AN(n4563), .B(n2777), .Y(N2791) );
  AOI21 U5456 ( .A0(n4682), .A1(n4683), .B0(n4684), .Y(n4563) );
  MX2 U5457 ( .A(n4685), .B(n4686), .S0(n4687), .Y(n4684) );
  NOR2 U5458 ( .A(in1_disp[29]), .B(n2679), .Y(n4686) );
  NOR2B U5459 ( .AN(n4688), .B(n4682), .Y(n4685) );
  NOR2B U5460 ( .AN(n4572), .B(n2780), .Y(N2790) );
  OAI211 U5461 ( .A0(in1_disp[29]), .A1(n4689), .B0(n4690), .C0(n4691), .Y(
        n4572) );
  INV U5462 ( .A(n4692), .Y(n4691) );
  MX2 U5463 ( .A(n4693), .B(n4694), .S0(n2619), .Y(n4690) );
  INV U5464 ( .A(n4688), .Y(n4694) );
  NOR2 U5465 ( .A(n4683), .B(n4589), .Y(n4693) );
  NOR2B U5466 ( .AN(n2679), .B(n4695), .Y(n4683) );
  INV U5467 ( .A(n4696), .Y(n4689) );
  NOR2 U5468 ( .A(n4581), .B(n2779), .Y(N2789) );
  NOR4 U5469 ( .A(n4682), .B(n4687), .C(n4697), .D(n4698), .Y(n4581) );
  NOR2B U5470 ( .AN(n2679), .B(n4699), .Y(n4698) );
  NOR2 U5471 ( .A(n2619), .B(in1_disp[29]), .Y(n4697) );
  NOR2B U5472 ( .AN(n4700), .B(n2778), .Y(N2788) );
  OAI31 U5473 ( .A0(n2679), .A1(n4695), .A2(n4589), .B0(n4590), .Y(n4700) );
  MX2 U5474 ( .A(n4701), .B(n4702), .S0(in1_disp[29]), .Y(n4590) );
  NOR3 U5475 ( .A(n2619), .B(n4692), .C(n4702), .Y(n4701) );
  NOR2 U5476 ( .A(n4696), .B(n4703), .Y(n4702) );
  NOR2B U5477 ( .AN(n2679), .B(in1_disp[30]), .Y(n4703) );
  NOR2 U5478 ( .A(n4594), .B(n2777), .Y(N2787) );
  NOR3B U5479 ( .AN(n4704), .B(n4692), .C(n4699), .Y(n4594) );
  NOR2 U5480 ( .A(in1_disp[30]), .B(n2679), .Y(n4692) );
  AOI22 U5481 ( .A0(in1_disp[30]), .A1(n2619), .B0(in1_disp[29]), .B1(n2678), 
        .Y(n4704) );
  NOR2 U5482 ( .A(n4598), .B(n2780), .Y(N2786) );
  NOR3 U5483 ( .A(n4682), .B(n4699), .C(n4705), .Y(n4598) );
  OAI2BB2 U5484 ( .B0(n2679), .B1(n4706), .A0N(n4687), .A1N(n4695), .Y(n4705)
         );
  NOR2B U5485 ( .AN(in1_disp[30]), .B(n2619), .Y(n4687) );
  NOR2 U5486 ( .A(in1_disp[30]), .B(n4695), .Y(n4706) );
  NOR2B U5487 ( .AN(n2619), .B(n4695), .Y(n4699) );
  NOR2B U5488 ( .AN(n2619), .B(in1_disp[30]), .Y(n4682) );
  NOR2 U5489 ( .A(n4600), .B(n2779), .Y(N2785) );
  NOR2 U5490 ( .A(enter), .B(n4961), .Y(n4161) );
  INV U5491 ( .A(data_type), .Y(n4961) );
  NOR2B U5492 ( .AN(n4707), .B(n4708), .Y(n4600) );
  AOI2BB1 U5493 ( .A0N(in1_disp[29]), .A1N(n4589), .B0(n2618), .Y(n4708) );
  MX2 U5494 ( .A(n4695), .B(n4709), .S0(in1_disp[30]), .Y(n4707) );
  NOR2 U5495 ( .A(n4688), .B(n4696), .Y(n4709) );
  NOR2 U5496 ( .A(n2619), .B(n2679), .Y(n4696) );
  NOR2B U5497 ( .AN(n2679), .B(in1_disp[29]), .Y(n4688) );
  OAI2BB2 U5498 ( .B0(n4710), .B1(n2770), .A0N(in2_disp[3]), .A1N(n2755), .Y(
        N2710) );
  NOR2 U5499 ( .A(in2_disp[3]), .B(n4711), .Y(n4710) );
  NOR2B U5500 ( .AN(n2559), .B(n2741), .Y(n4711) );
  OAI2BB2 U5501 ( .B0(n2754), .B1(n2616), .A0N(n2559), .A1N(n2657), .Y(N2709)
         );
  OAI2BB2 U5502 ( .B0(n2754), .B1(n4715), .A0N(n2559), .A1N(n2650), .Y(N2708)
         );
  INV U5503 ( .A(in2_disp[1]), .Y(n4715) );
  OAI2BB2 U5504 ( .B0(n4716), .B1(n2770), .A0N(n2615), .A1N(n2755), .Y(N2707)
         );
  NOR2 U5505 ( .A(n2615), .B(n4717), .Y(n4716) );
  NOR2B U5506 ( .AN(n2559), .B(n2731), .Y(n4717) );
  NOR3B U5507 ( .AN(input2_cnt[1]), .B(n4719), .C(n3447), .Y(n3449) );
  OAI2BB2 U5508 ( .B0(n4720), .B1(n2770), .A0N(in2_disp[7]), .A1N(n2755), .Y(
        N2706) );
  NOR2 U5509 ( .A(in2_disp[7]), .B(n4721), .Y(n4720) );
  NOR2B U5510 ( .AN(n4722), .B(n2741), .Y(n4721) );
  OAI2BB2 U5511 ( .B0(n2754), .B1(n2612), .A0N(n2657), .A1N(n4722), .Y(N2705)
         );
  OAI2BB2 U5512 ( .B0(n2754), .B1(n4723), .A0N(n2650), .A1N(n4722), .Y(N2704)
         );
  INV U5513 ( .A(in2_disp[5]), .Y(n4723) );
  OAI2BB2 U5514 ( .B0(n4724), .B1(n2770), .A0N(n2611), .A1N(n2755), .Y(N2703)
         );
  NOR2 U5515 ( .A(n2611), .B(n4725), .Y(n4724) );
  NOR2B U5516 ( .AN(n4722), .B(n2731), .Y(n4725) );
  NOR2B U5517 ( .AN(n4726), .B(n4719), .Y(n4722) );
  OAI2BB2 U5518 ( .B0(n4727), .B1(n2770), .A0N(in2_disp[11]), .A1N(n2755), .Y(
        N2702) );
  NOR2 U5519 ( .A(in2_disp[11]), .B(n4728), .Y(n4727) );
  NOR2B U5520 ( .AN(n4729), .B(n2741), .Y(n4728) );
  OAI2BB2 U5521 ( .B0(n2754), .B1(n4247), .A0N(n2657), .A1N(n4729), .Y(N2701)
         );
  INV U5522 ( .A(in2_disp[10]), .Y(n4247) );
  OAI2BB2 U5523 ( .B0(n2754), .B1(n4242), .A0N(n2650), .A1N(n4729), .Y(N2700)
         );
  INV U5524 ( .A(in2_disp[9]), .Y(n4242) );
  OAI2BB2 U5525 ( .B0(n4730), .B1(n2770), .A0N(in2_disp[8]), .A1N(n2755), .Y(
        N2699) );
  NOR2 U5526 ( .A(in2_disp[8]), .B(n4731), .Y(n4730) );
  NOR2B U5527 ( .AN(n4729), .B(n2731), .Y(n4731) );
  NOR3 U5528 ( .A(input2_cnt[1]), .B(n4719), .C(n3447), .Y(n4729) );
  OAI2BB2 U5529 ( .B0(n4732), .B1(n2770), .A0N(in2_disp[15]), .A1N(n2755), .Y(
        N2698) );
  NOR2 U5530 ( .A(in2_disp[15]), .B(n4733), .Y(n4732) );
  NOR2B U5531 ( .AN(n4734), .B(n2741), .Y(n4733) );
  OAI2BB2 U5532 ( .B0(n2754), .B1(n2608), .A0N(n2657), .A1N(n4734), .Y(N2697)
         );
  OAI2BB2 U5533 ( .B0(n2754), .B1(n4735), .A0N(n2650), .A1N(n4734), .Y(N2696)
         );
  INV U5534 ( .A(in2_disp[13]), .Y(n4735) );
  OAI2BB2 U5535 ( .B0(n4736), .B1(n2770), .A0N(n2607), .A1N(n2755), .Y(N2695)
         );
  NOR2 U5536 ( .A(n2607), .B(n4737), .Y(n4736) );
  NOR2B U5537 ( .AN(n4734), .B(n2731), .Y(n4737) );
  NOR3 U5538 ( .A(input2_cnt[0]), .B(input2_cnt[1]), .C(n4719), .Y(n4734) );
  OAI2BB2 U5539 ( .B0(n4738), .B1(n2770), .A0N(n2605), .A1N(n2755), .Y(N2694)
         );
  NOR2 U5540 ( .A(n2605), .B(n4739), .Y(n4738) );
  NOR2B U5541 ( .AN(n4740), .B(n2741), .Y(n4739) );
  OAI2BB2 U5542 ( .B0(n2754), .B1(n4171), .A0N(n2657), .A1N(n4740), .Y(N2693)
         );
  INV U5543 ( .A(in2_disp[18]), .Y(n4171) );
  OAI2BB2 U5544 ( .B0(n2754), .B1(n4335), .A0N(n2650), .A1N(n4740), .Y(N2692)
         );
  INV U5545 ( .A(in2_disp[17]), .Y(n4335) );
  OAI2BB2 U5546 ( .B0(n4741), .B1(n2770), .A0N(n2677), .A1N(n2755), .Y(N2691)
         );
  NOR2 U5547 ( .A(n2677), .B(n4742), .Y(n4741) );
  NOR2B U5548 ( .AN(n4740), .B(n2731), .Y(n4742) );
  NOR3B U5549 ( .AN(input2_cnt[1]), .B(input2_cnt[2]), .C(n3447), .Y(n4740) );
  OAI2BB2 U5550 ( .B0(n4743), .B1(n2770), .A0N(n2603), .A1N(n2755), .Y(N2690)
         );
  NOR2 U5551 ( .A(n2603), .B(n4744), .Y(n4743) );
  NOR2B U5552 ( .AN(n4745), .B(n2741), .Y(n4744) );
  OAI2BB2 U5553 ( .B0(n2754), .B1(n4217), .A0N(n2657), .A1N(n4745), .Y(N2689)
         );
  INV U5554 ( .A(in2_disp[22]), .Y(n4217) );
  OAI2BB2 U5555 ( .B0(n2754), .B1(n4363), .A0N(n2650), .A1N(n4745), .Y(N2688)
         );
  INV U5556 ( .A(in2_disp[21]), .Y(n4363) );
  OAI2BB2 U5557 ( .B0(n4746), .B1(n2770), .A0N(n2683), .A1N(n2755), .Y(N2687)
         );
  NOR2 U5558 ( .A(n2683), .B(n4747), .Y(n4746) );
  NOR2B U5559 ( .AN(n4745), .B(n2731), .Y(n4747) );
  NOR2B U5560 ( .AN(n4726), .B(input2_cnt[2]), .Y(n4745) );
  NOR2B U5561 ( .AN(input2_cnt[1]), .B(input2_cnt[0]), .Y(n4726) );
  OAI2BB2 U5562 ( .B0(n4748), .B1(n2770), .A0N(n2601), .A1N(n2755), .Y(N2686)
         );
  NOR2 U5563 ( .A(n2601), .B(n4749), .Y(n4748) );
  NOR2B U5564 ( .AN(n4750), .B(n2741), .Y(n4749) );
  OAI2BB2 U5565 ( .B0(n2754), .B1(n4390), .A0N(n2657), .A1N(n4750), .Y(N2685)
         );
  INV U5566 ( .A(in2_disp[26]), .Y(n4390) );
  OAI2BB2 U5567 ( .B0(n2754), .B1(n4751), .A0N(n2650), .A1N(n4750), .Y(N2684)
         );
  INV U5568 ( .A(in2_disp[25]), .Y(n4751) );
  OAI2BB2 U5569 ( .B0(n4752), .B1(n2770), .A0N(in2_disp[24]), .A1N(n2755), .Y(
        N2683) );
  NOR2 U5570 ( .A(in2_disp[24]), .B(n4753), .Y(n4752) );
  NOR2B U5571 ( .AN(n4750), .B(n2731), .Y(n4753) );
  NOR2B U5572 ( .AN(n4754), .B(n3447), .Y(n4750) );
  INV U5573 ( .A(input2_cnt[0]), .Y(n3447) );
  OAI2BB2 U5574 ( .B0(n4755), .B1(n2770), .A0N(n2599), .A1N(n2755), .Y(N2682)
         );
  NOR2 U5575 ( .A(n2599), .B(n4756), .Y(n4755) );
  NOR2B U5576 ( .AN(n4757), .B(n2741), .Y(n4756) );
  NOR4BB U5577 ( .AN(n4758), .BN(n4759), .C(n4760), .D(n4761), .Y(n4712) );
  AOI21 U5578 ( .A0(n4762), .A1(n4763), .B0(n4764), .Y(n4759) );
  OAI2BB2 U5579 ( .B0(n2754), .B1(n4307), .A0N(n2657), .A1N(n4757), .Y(N2681)
         );
  AOI31 U5580 ( .A0(n4765), .A1(n4766), .A2(n4767), .B0(n2770), .Y(n4714) );
  AOI211 U5581 ( .A0(n4762), .A1(n4768), .B0(n4769), .C0(n4764), .Y(n4765) );
  NOR2B U5582 ( .AN(n4770), .B(n4771), .Y(n4764) );
  INV U5583 ( .A(n4772), .Y(n4762) );
  INV U5584 ( .A(in2_disp[30]), .Y(n4307) );
  OAI2BB2 U5585 ( .B0(n2754), .B1(n4413), .A0N(n2650), .A1N(n4757), .Y(N2680)
         );
  NOR4B U5586 ( .AN(n4758), .B(n4774), .C(n4775), .D(n4776), .Y(n4773) );
  OAI2BB1 U5587 ( .A0N(n4777), .A1N(n4768), .B0(n4767), .Y(n4776) );
  NAND2 U5588 ( .A(n4777), .B(n4763), .Y(n4767) );
  INV U5589 ( .A(n4778), .Y(n4768) );
  NOR4 U5590 ( .A(n4779), .B(n4780), .C(n4769), .D(n4781), .Y(n4758) );
  NOR2B U5591 ( .AN(n4782), .B(n4783), .Y(n4781) );
  NOR2B U5592 ( .AN(n4770), .B(n4783), .Y(n4769) );
  INV U5593 ( .A(in2_disp[29]), .Y(n4413) );
  NOR2B U5594 ( .AN(ce), .B(n2769), .Y(n4713) );
  OAI2BB2 U5595 ( .B0(n4784), .B1(n2770), .A0N(n2681), .A1N(n2755), .Y(N2679)
         );
  OAI211 U5596 ( .A0(data_type), .A1(n4719), .B0(n4785), .C0(n4786), .Y(n3446)
         );
  AOI2BB2 U5597 ( .B0(n4787), .B1(n4788), .A0N(in2_row_reg[3]), .A1N(n4778), 
        .Y(n4785) );
  INV U5598 ( .A(in2_col_reg[1]), .Y(n4788) );
  INV U5599 ( .A(n4783), .Y(n4787) );
  INV U5600 ( .A(input2_cnt[2]), .Y(n4719) );
  NOR2 U5601 ( .A(n2681), .B(n4789), .Y(n4784) );
  NOR2B U5602 ( .AN(n4757), .B(n2731), .Y(n4789) );
  NOR4BB U5603 ( .AN(n4766), .BN(n4790), .C(n4780), .D(n4761), .Y(n4718) );
  NOR2B U5604 ( .AN(n4782), .B(n4771), .Y(n4761) );
  NOR2B U5605 ( .AN(n4782), .B(n4772), .Y(n4780) );
  NOR3 U5606 ( .A(in2_row_reg[3]), .B(in2_row_reg[0]), .C(in2_row_reg[2]), .Y(
        n4782) );
  AOI2BB1 U5607 ( .A0N(n4771), .A1N(n4778), .B0(n4774), .Y(n4790) );
  NOR2 U5608 ( .A(n4778), .B(n4783), .Y(n4774) );
  NAND2B U5609 ( .AN(in2_row_reg[0]), .B(n4791), .Y(n4778) );
  NOR4 U5610 ( .A(n4779), .B(n4760), .C(n4775), .D(n4792), .Y(n4766) );
  NOR2B U5611 ( .AN(n4763), .B(n4771), .Y(n4792) );
  OR3 U5612 ( .A(in2_col_reg[1]), .B(in2_col_reg[0]), .C(in2_col_reg[2]), .Y(
        n4771) );
  NOR2B U5613 ( .AN(n4763), .B(n4783), .Y(n4775) );
  NAND2B U5614 ( .AN(in2_col_reg[0]), .B(n4793), .Y(n4783) );
  NOR3 U5615 ( .A(in2_row_reg[3]), .B(in2_row_reg[0]), .C(in2_row_reg[1]), .Y(
        n4763) );
  NOR2B U5616 ( .AN(n4777), .B(n4794), .Y(n4760) );
  INV U5617 ( .A(n4770), .Y(n4794) );
  NOR3 U5618 ( .A(in2_col_reg[1]), .B(in2_col_reg[0]), .C(in2_col_reg[3]), .Y(
        n4777) );
  NOR2B U5619 ( .AN(n4770), .B(n4772), .Y(n4779) );
  NAND2B U5620 ( .AN(in2_col_reg[1]), .B(n4793), .Y(n4772) );
  NOR2 U5621 ( .A(in2_col_reg[3]), .B(in2_col_reg[2]), .Y(n4793) );
  NOR2B U5622 ( .AN(n4791), .B(in2_row_reg[3]), .Y(n4770) );
  NOR2 U5623 ( .A(in2_row_reg[2]), .B(in2_row_reg[1]), .Y(n4791) );
  NOR2B U5624 ( .AN(n4754), .B(input2_cnt[0]), .Y(n4757) );
  NOR2 U5625 ( .A(input2_cnt[2]), .B(input2_cnt[1]), .Y(n4754) );
  OAI2BB2 U5626 ( .B0(n4795), .B1(n2772), .A0N(in1_disp[3]), .A1N(n2744), .Y(
        N1451) );
  NOR2 U5627 ( .A(in1_disp[3]), .B(n4796), .Y(n4795) );
  NOR2B U5628 ( .AN(n2561), .B(n2733), .Y(n4796) );
  OAI2BB2 U5629 ( .B0(n2743), .B1(n2636), .A0N(n2561), .A1N(n2659), .Y(N1450)
         );
  OAI2BB2 U5630 ( .B0(n2743), .B1(n4800), .A0N(n2561), .A1N(n2651), .Y(N1449)
         );
  INV U5631 ( .A(in1_disp[1]), .Y(n4800) );
  OAI2BB2 U5632 ( .B0(n4801), .B1(n2772), .A0N(n2635), .A1N(n2744), .Y(N1448)
         );
  NOR2 U5633 ( .A(n2635), .B(n4802), .Y(n4801) );
  NOR2B U5634 ( .AN(n2561), .B(n2727), .Y(n4802) );
  NOR3B U5635 ( .AN(input1_cnt[1]), .B(n4804), .C(n3437), .Y(n3439) );
  OAI2BB2 U5636 ( .B0(n4805), .B1(n2772), .A0N(in1_disp[7]), .A1N(n2744), .Y(
        N1447) );
  NOR2 U5637 ( .A(in1_disp[7]), .B(n4806), .Y(n4805) );
  NOR2B U5638 ( .AN(n4807), .B(n2733), .Y(n4806) );
  OAI2BB2 U5639 ( .B0(n2743), .B1(n2632), .A0N(n2659), .A1N(n4807), .Y(N1446)
         );
  OAI2BB2 U5640 ( .B0(n2743), .B1(n4808), .A0N(n2651), .A1N(n4807), .Y(N1445)
         );
  INV U5641 ( .A(in1_disp[5]), .Y(n4808) );
  OAI2BB2 U5642 ( .B0(n4809), .B1(n2772), .A0N(n2631), .A1N(n2744), .Y(N1444)
         );
  NOR2 U5643 ( .A(n2631), .B(n4810), .Y(n4809) );
  NOR2B U5644 ( .AN(n4807), .B(n2727), .Y(n4810) );
  NOR2B U5645 ( .AN(n4811), .B(n4804), .Y(n4807) );
  OAI2BB2 U5646 ( .B0(n4812), .B1(n2772), .A0N(in1_disp[11]), .A1N(n2744), .Y(
        N1443) );
  NOR2 U5647 ( .A(in1_disp[11]), .B(n4813), .Y(n4812) );
  NOR2B U5648 ( .AN(n4814), .B(n2733), .Y(n4813) );
  OAI2BB2 U5649 ( .B0(n2743), .B1(n4529), .A0N(n2659), .A1N(n4814), .Y(N1442)
         );
  INV U5650 ( .A(in1_disp[10]), .Y(n4529) );
  OAI2BB2 U5651 ( .B0(n2743), .B1(n4524), .A0N(n2651), .A1N(n4814), .Y(N1441)
         );
  INV U5652 ( .A(in1_disp[9]), .Y(n4524) );
  OAI2BB2 U5653 ( .B0(n4815), .B1(n2772), .A0N(in1_disp[8]), .A1N(n2744), .Y(
        N1440) );
  NOR2 U5654 ( .A(in1_disp[8]), .B(n4816), .Y(n4815) );
  NOR2B U5655 ( .AN(n4814), .B(n2727), .Y(n4816) );
  NOR3 U5656 ( .A(input1_cnt[1]), .B(n4804), .C(n3437), .Y(n4814) );
  OAI2BB2 U5657 ( .B0(n4817), .B1(n2772), .A0N(in1_disp[15]), .A1N(n2744), .Y(
        N1439) );
  NOR2 U5658 ( .A(in1_disp[15]), .B(n4818), .Y(n4817) );
  NOR2B U5659 ( .AN(n4819), .B(n2733), .Y(n4818) );
  OAI2BB2 U5660 ( .B0(n2743), .B1(n2628), .A0N(n2659), .A1N(n4819), .Y(N1438)
         );
  OAI2BB2 U5661 ( .B0(n2743), .B1(n4820), .A0N(n2651), .A1N(n4819), .Y(N1437)
         );
  INV U5662 ( .A(in1_disp[13]), .Y(n4820) );
  OAI2BB2 U5663 ( .B0(n4821), .B1(n2772), .A0N(n2627), .A1N(n2744), .Y(N1436)
         );
  NOR2 U5664 ( .A(n2627), .B(n4822), .Y(n4821) );
  NOR2B U5665 ( .AN(n4819), .B(n2727), .Y(n4822) );
  NOR3 U5666 ( .A(input1_cnt[0]), .B(input1_cnt[1]), .C(n4804), .Y(n4819) );
  OAI2BB2 U5667 ( .B0(n4823), .B1(n2772), .A0N(n2625), .A1N(n2744), .Y(N1435)
         );
  NOR2 U5668 ( .A(n2625), .B(n4824), .Y(n4823) );
  NOR2B U5669 ( .AN(n4825), .B(n2733), .Y(n4824) );
  OAI2BB2 U5670 ( .B0(n2743), .B1(n4457), .A0N(n2659), .A1N(n4825), .Y(N1434)
         );
  INV U5671 ( .A(in1_disp[18]), .Y(n4457) );
  OAI2BB2 U5672 ( .B0(n2743), .B1(n4617), .A0N(n2651), .A1N(n4825), .Y(N1433)
         );
  INV U5673 ( .A(in1_disp[17]), .Y(n4617) );
  OAI2BB2 U5674 ( .B0(n4826), .B1(n2772), .A0N(n2675), .A1N(n2744), .Y(N1432)
         );
  NOR2 U5675 ( .A(n2675), .B(n4827), .Y(n4826) );
  NOR2B U5676 ( .AN(n4825), .B(n2727), .Y(n4827) );
  NOR3B U5677 ( .AN(input1_cnt[1]), .B(input1_cnt[2]), .C(n3437), .Y(n4825) );
  OAI2BB2 U5678 ( .B0(n4828), .B1(n2772), .A0N(n2623), .A1N(n2744), .Y(N1431)
         );
  NOR2 U5679 ( .A(n2623), .B(n4829), .Y(n4828) );
  NOR2B U5680 ( .AN(n4830), .B(n2733), .Y(n4829) );
  OAI2BB2 U5681 ( .B0(n2743), .B1(n4501), .A0N(n2659), .A1N(n4830), .Y(N1430)
         );
  INV U5682 ( .A(in1_disp[22]), .Y(n4501) );
  OAI2BB2 U5683 ( .B0(n2743), .B1(n4645), .A0N(n2651), .A1N(n4830), .Y(N1429)
         );
  INV U5684 ( .A(in1_disp[21]), .Y(n4645) );
  OAI2BB2 U5685 ( .B0(n4831), .B1(n2772), .A0N(n2673), .A1N(n2744), .Y(N1428)
         );
  NOR2 U5686 ( .A(n2673), .B(n4832), .Y(n4831) );
  NOR2B U5687 ( .AN(n4830), .B(n2727), .Y(n4832) );
  NOR2B U5688 ( .AN(n4811), .B(input1_cnt[2]), .Y(n4830) );
  NOR2B U5689 ( .AN(input1_cnt[1]), .B(input1_cnt[0]), .Y(n4811) );
  OAI2BB2 U5690 ( .B0(n4833), .B1(n2772), .A0N(n2621), .A1N(n2744), .Y(N1427)
         );
  NOR2 U5691 ( .A(n2621), .B(n4834), .Y(n4833) );
  NOR2B U5692 ( .AN(n4835), .B(n2733), .Y(n4834) );
  OAI2BB2 U5693 ( .B0(n2743), .B1(n4672), .A0N(n2659), .A1N(n4835), .Y(N1426)
         );
  INV U5694 ( .A(in1_disp[26]), .Y(n4672) );
  OAI2BB2 U5695 ( .B0(n2743), .B1(n4836), .A0N(n2651), .A1N(n4835), .Y(N1425)
         );
  INV U5696 ( .A(in1_disp[25]), .Y(n4836) );
  OAI2BB2 U5697 ( .B0(n4837), .B1(n2772), .A0N(in1_disp[24]), .A1N(n2744), .Y(
        N1424) );
  NOR2 U5698 ( .A(in1_disp[24]), .B(n4838), .Y(n4837) );
  NOR2B U5699 ( .AN(n4835), .B(n2727), .Y(n4838) );
  NOR2B U5700 ( .AN(n4839), .B(n3437), .Y(n4835) );
  INV U5701 ( .A(input1_cnt[0]), .Y(n3437) );
  OAI2BB2 U5702 ( .B0(n4840), .B1(n2772), .A0N(n2619), .A1N(n2744), .Y(N1423)
         );
  NOR2 U5703 ( .A(n2619), .B(n4841), .Y(n4840) );
  NOR2B U5704 ( .AN(n4842), .B(n2733), .Y(n4841) );
  NOR4BB U5705 ( .AN(n4843), .BN(n4844), .C(n4845), .D(n4846), .Y(n4797) );
  AOI21 U5706 ( .A0(n4847), .A1(n4848), .B0(n4849), .Y(n4844) );
  OAI2BB2 U5707 ( .B0(n2743), .B1(n4589), .A0N(n2659), .A1N(n4842), .Y(N1422)
         );
  AOI31 U5708 ( .A0(n4850), .A1(n4851), .A2(n4852), .B0(n2772), .Y(n4799) );
  AOI211 U5709 ( .A0(n4847), .A1(n4853), .B0(n4854), .C0(n4849), .Y(n4850) );
  NOR2B U5710 ( .AN(n4855), .B(n4856), .Y(n4849) );
  INV U5711 ( .A(n4857), .Y(n4847) );
  INV U5712 ( .A(in1_disp[30]), .Y(n4589) );
  OAI2BB2 U5713 ( .B0(n2743), .B1(n4695), .A0N(n2651), .A1N(n4842), .Y(N1421)
         );
  NOR4B U5714 ( .AN(n4843), .B(n4859), .C(n4860), .D(n4861), .Y(n4858) );
  OAI2BB1 U5715 ( .A0N(n4862), .A1N(n4853), .B0(n4852), .Y(n4861) );
  NAND2 U5716 ( .A(n4862), .B(n4848), .Y(n4852) );
  INV U5717 ( .A(n4863), .Y(n4853) );
  NOR4 U5718 ( .A(n4864), .B(n4865), .C(n4854), .D(n4866), .Y(n4843) );
  NOR2B U5719 ( .AN(n4867), .B(n4868), .Y(n4866) );
  NOR2B U5720 ( .AN(n4855), .B(n4868), .Y(n4854) );
  INV U5721 ( .A(in1_disp[29]), .Y(n4695) );
  NOR2B U5722 ( .AN(ce), .B(n2771), .Y(n4798) );
  OAI2BB2 U5723 ( .B0(n4869), .B1(n2772), .A0N(n2679), .A1N(n2744), .Y(N1420)
         );
  OAI211 U5724 ( .A0(data_type), .A1(n4804), .B0(n4870), .C0(n4871), .Y(n3436)
         );
  AOI2BB2 U5725 ( .B0(n4872), .B1(n4873), .A0N(in1_row_reg[3]), .A1N(n4863), 
        .Y(n4870) );
  INV U5726 ( .A(in1_col_reg[1]), .Y(n4873) );
  INV U5727 ( .A(n4868), .Y(n4872) );
  INV U5728 ( .A(input1_cnt[2]), .Y(n4804) );
  NOR2 U5729 ( .A(n2679), .B(n4874), .Y(n4869) );
  NOR2B U5730 ( .AN(n4842), .B(n2727), .Y(n4874) );
  NOR4BB U5731 ( .AN(n4851), .BN(n4875), .C(n4865), .D(n4846), .Y(n4803) );
  NOR2B U5732 ( .AN(n4867), .B(n4856), .Y(n4846) );
  NOR2B U5733 ( .AN(n4867), .B(n4857), .Y(n4865) );
  NOR3 U5734 ( .A(in1_row_reg[3]), .B(in1_row_reg[0]), .C(in1_row_reg[2]), .Y(
        n4867) );
  AOI2BB1 U5735 ( .A0N(n4856), .A1N(n4863), .B0(n4859), .Y(n4875) );
  NOR2 U5736 ( .A(n4863), .B(n4868), .Y(n4859) );
  NAND2B U5737 ( .AN(in1_row_reg[0]), .B(n4876), .Y(n4863) );
  NOR4 U5738 ( .A(n4864), .B(n4845), .C(n4860), .D(n4877), .Y(n4851) );
  NOR2B U5739 ( .AN(n4848), .B(n4856), .Y(n4877) );
  OR3 U5740 ( .A(in1_col_reg[1]), .B(in1_col_reg[0]), .C(in1_col_reg[2]), .Y(
        n4856) );
  NOR2B U5741 ( .AN(n4848), .B(n4868), .Y(n4860) );
  NAND2B U5742 ( .AN(in1_col_reg[0]), .B(n4878), .Y(n4868) );
  NOR3 U5743 ( .A(in1_row_reg[3]), .B(in1_row_reg[0]), .C(in1_row_reg[1]), .Y(
        n4848) );
  NOR2B U5744 ( .AN(n4862), .B(n4879), .Y(n4845) );
  INV U5745 ( .A(n4855), .Y(n4879) );
  NOR3 U5746 ( .A(in1_col_reg[1]), .B(in1_col_reg[0]), .C(in1_col_reg[3]), .Y(
        n4862) );
  NOR2B U5747 ( .AN(n4855), .B(n4857), .Y(n4864) );
  NAND2B U5748 ( .AN(in1_col_reg[1]), .B(n4878), .Y(n4857) );
  NOR2 U5749 ( .A(in1_col_reg[3]), .B(in1_col_reg[2]), .Y(n4878) );
  NOR2B U5750 ( .AN(n4876), .B(in1_row_reg[3]), .Y(n4855) );
  NOR2 U5751 ( .A(in1_row_reg[2]), .B(in1_row_reg[1]), .Y(n4876) );
  NOR2B U5752 ( .AN(n4839), .B(input1_cnt[0]), .Y(n4842) );
  NOR2 U5753 ( .A(input1_cnt[2]), .B(input1_cnt[1]), .Y(n4839) );
endmodule

